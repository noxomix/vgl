module vgl

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="AttribMask" type="bitmask" |>
pub const (
	gl_current_bit          = int(0x00000001)
	gl_point_bit            = int(0x00000002)
	gl_line_bit             = int(0x00000004)
	gl_polygon_bit          = int(0x00000008)
	gl_polygon_stipple_bit  = int(0x00000010)
	gl_pixel_mode_bit       = int(0x00000020)
	gl_lighting_bit         = int(0x00000040)
	gl_fog_bit              = int(0x00000080)
	gl_depth_buffer_bit     = int(0x00000100)
	gl_accum_buffer_bit     = int(0x00000200)
	gl_stencil_buffer_bit   = int(0x00000400)
	gl_viewport_bit         = int(0x00000800)
	gl_transform_bit        = int(0x00001000)
	gl_enable_bit           = int(0x00002000)
	gl_color_buffer_bit     = int(0x00004000)
	gl_hint_bit             = int(0x00008000)
	gl_eval_bit             = int(0x00010000)
	gl_list_bit             = int(0x00020000)
	gl_texture_bit          = int(0x00040000)
	gl_scissor_bit          = int(0x00080000)
	gl_multisample_bit      = int(0x20000000)
	gl_multisample_bit_arb  = int(0x20000000)
	gl_multisample_bit_ext  = int(0x20000000)
	gl_multisample_bit_3dfx = int(0x20000000)
	gl_all_attrib_bits      = int(0xFFFFFFFF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="BufferStorageMask" type="bitmask" comment="GL_MAP_{COHERENT,PERSISTENT,READ,WRITE}_{BIT,BIT_EXT} also lie in this namespace" |>
pub const (
	gl_dynamic_storage_bit           = int(0x0100)
	gl_dynamic_storage_bit_ext       = int(0x0100)
	gl_client_storage_bit            = int(0x0200)
	gl_client_storage_bit_ext        = int(0x0200)
	gl_sparse_storage_bit_arb        = int(0x0400)
	gl_lgpu_separate_storage_bit_nvx = int(0x0800)
	gl_per_gpu_storage_bit_nv        = int(0x0800)
	gl_external_storage_bit_nvx      = int(0x2000)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="ClearBufferMask" type="bitmask" comment="GL_{DEPTH,ACCUM,STENCIL,COLOR}_BUFFER_BIT also lie in this namespace" |>
pub const (
	gl_coverage_buffer_bit_nv = int(0x00008000)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="ClientAttribMask" type="bitmask" |>
pub const (
	gl_client_pixel_store_bit  = int(0x00000001)
	gl_client_vertex_array_bit = int(0x00000002)
	gl_client_all_attrib_bits  = int(0xFFFFFFFF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="ContextFlagMask" type="bitmask" comment="Should be shared with WGL/GLX, but aren't since the FORWARD_COMPATIBLE and DEBUG values are swapped vs. WGL/GLX." |>
pub const (
	gl_context_flag_forward_compatible_bit    = int(0x00000001)
	gl_context_flag_debug_bit                 = int(0x00000002)
	gl_context_flag_debug_bit_khr             = int(0x00000002)
	gl_context_flag_robust_access_bit         = int(0x00000004)
	gl_context_flag_robust_access_bit_arb     = int(0x00000004)
	gl_context_flag_no_error_bit              = int(0x00000008)
	gl_context_flag_no_error_bit_khr          = int(0x00000008)
	gl_context_flag_protected_content_bit_ext = int(0x00000010)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="ContextProfileMask" type="bitmask" |>
pub const (
	gl_context_core_profile_bit          = int(0x00000001)
	gl_context_compatibility_profile_bit = int(0x00000002)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="MapBufferAccessMask" type="bitmask" |>
pub const (
	gl_map_read_bit                  = int(0x0001)
	gl_map_read_bit_ext              = int(0x0001)
	gl_map_write_bit                 = int(0x0002)
	gl_map_write_bit_ext             = int(0x0002)
	gl_map_invalidate_range_bit      = int(0x0004)
	gl_map_invalidate_range_bit_ext  = int(0x0004)
	gl_map_invalidate_buffer_bit     = int(0x0008)
	gl_map_invalidate_buffer_bit_ext = int(0x0008)
	gl_map_flush_explicit_bit        = int(0x0010)
	gl_map_flush_explicit_bit_ext    = int(0x0010)
	gl_map_unsynchronized_bit        = int(0x0020)
	gl_map_unsynchronized_bit_ext    = int(0x0020)
	gl_map_persistent_bit            = int(0x0040)
	gl_map_persistent_bit_ext        = int(0x0040)
	gl_map_coherent_bit              = int(0x0080)
	gl_map_coherent_bit_ext          = int(0x0080)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="MemoryBarrierMask" type="bitmask" |>
pub const (
	gl_vertex_attrib_array_barrier_bit      = int(0x00000001)
	gl_vertex_attrib_array_barrier_bit_ext  = int(0x00000001)
	gl_element_array_barrier_bit            = int(0x00000002)
	gl_element_array_barrier_bit_ext        = int(0x00000002)
	gl_uniform_barrier_bit                  = int(0x00000004)
	gl_uniform_barrier_bit_ext              = int(0x00000004)
	gl_texture_fetch_barrier_bit            = int(0x00000008)
	gl_texture_fetch_barrier_bit_ext        = int(0x00000008)
	gl_shader_global_access_barrier_bit_nv  = int(0x00000010)
	gl_shader_image_access_barrier_bit      = int(0x00000020)
	gl_shader_image_access_barrier_bit_ext  = int(0x00000020)
	gl_command_barrier_bit                  = int(0x00000040)
	gl_command_barrier_bit_ext              = int(0x00000040)
	gl_pixel_buffer_barrier_bit             = int(0x00000080)
	gl_pixel_buffer_barrier_bit_ext         = int(0x00000080)
	gl_texture_update_barrier_bit           = int(0x00000100)
	gl_texture_update_barrier_bit_ext       = int(0x00000100)
	gl_buffer_update_barrier_bit            = int(0x00000200)
	gl_buffer_update_barrier_bit_ext        = int(0x00000200)
	gl_framebuffer_barrier_bit              = int(0x00000400)
	gl_framebuffer_barrier_bit_ext          = int(0x00000400)
	gl_transform_feedback_barrier_bit       = int(0x00000800)
	gl_transform_feedback_barrier_bit_ext   = int(0x00000800)
	gl_atomic_counter_barrier_bit           = int(0x00001000)
	gl_atomic_counter_barrier_bit_ext       = int(0x00001000)
	gl_shader_storage_barrier_bit           = int(0x00002000)
	gl_client_mapped_buffer_barrier_bit     = int(0x00004000)
	gl_client_mapped_buffer_barrier_bit_ext = int(0x00004000)
	gl_query_buffer_barrier_bit             = int(0x00008000)
	gl_all_barrier_bits                     = int(0xFFFFFFFF)
	gl_all_barrier_bits_ext                 = int(0xFFFFFFFF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="OcclusionQueryEventMaskAMD" type="bitmask" |>
pub const (
	gl_query_depth_pass_event_bit_amd        = int(0x00000001)
	gl_query_depth_fail_event_bit_amd        = int(0x00000002)
	gl_query_stencil_fail_event_bit_amd      = int(0x00000004)
	gl_query_depth_bounds_fail_event_bit_amd = int(0x00000008)
	gl_query_all_event_bits_amd              = int(0xFFFFFFFF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="SyncObjectMask" type="bitmask" |>
pub const (
	gl_sync_flush_commands_bit       = int(0x00000001)
	gl_sync_flush_commands_bit_apple = int(0x00000001)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="UseProgramStageMask" type="bitmask" |>
pub const (
	gl_vertex_shader_bit              = int(0x00000001)
	gl_vertex_shader_bit_ext          = int(0x00000001)
	gl_fragment_shader_bit            = int(0x00000002)
	gl_fragment_shader_bit_ext        = int(0x00000002)
	gl_geometry_shader_bit            = int(0x00000004)
	gl_geometry_shader_bit_ext        = int(0x00000004)
	gl_geometry_shader_bit_oes        = int(0x00000004)
	gl_tess_control_shader_bit        = int(0x00000008)
	gl_tess_control_shader_bit_ext    = int(0x00000008)
	gl_tess_control_shader_bit_oes    = int(0x00000008)
	gl_tess_evaluation_shader_bit     = int(0x00000010)
	gl_tess_evaluation_shader_bit_ext = int(0x00000010)
	gl_tess_evaluation_shader_bit_oes = int(0x00000010)
	gl_compute_shader_bit             = int(0x00000020)
	gl_mesh_shader_bit_nv             = int(0x00000040)
	gl_task_shader_bit_nv             = int(0x00000080)
	gl_all_shader_bits                = int(0xFFFFFFFF)
	gl_all_shader_bits_ext            = int(0xFFFFFFFF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="SubgroupSupportedFeatures" type="bitmask" |>
pub const (
	gl_subgroup_feature_basic_bit_khr            = int(0x00000001)
	gl_subgroup_feature_vote_bit_khr             = int(0x00000002)
	gl_subgroup_feature_arithmetic_bit_khr       = int(0x00000004)
	gl_subgroup_feature_ballot_bit_khr           = int(0x00000008)
	gl_subgroup_feature_shuffle_bit_khr          = int(0x00000010)
	gl_subgroup_feature_shuffle_relative_bit_khr = int(0x00000020)
	gl_subgroup_feature_clustered_bit_khr        = int(0x00000040)
	gl_subgroup_feature_quad_bit_khr             = int(0x00000080)
	gl_subgroup_feature_partitioned_bit_nv       = int(0x00000100)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="TextureStorageMaskAMD" type="bitmask" |>
pub const (
	gl_texture_storage_sparse_bit_amd = int(0x00000001)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="FragmentShaderDestMaskATI" type="bitmask" |>
pub const (
	gl_red_bit_ati   = int(0x00000001)
	gl_green_bit_ati = int(0x00000002)
	gl_blue_bit_ati  = int(0x00000004)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="FragmentShaderDestModMaskATI" type="bitmask" |>
pub const (
	gl_2x_bit_ati       = int(0x00000001)
	gl_4x_bit_ati       = int(0x00000002)
	gl_8x_bit_ati       = int(0x00000004)
	gl_half_bit_ati     = int(0x00000008)
	gl_quarter_bit_ati  = int(0x00000010)
	gl_eighth_bit_ati   = int(0x00000020)
	gl_saturate_bit_ati = int(0x00000040)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="FragmentShaderColorModMaskATI" type="bitmask" |>
pub const (
	gl_comp_bit_ati   = int(0x00000002)
	gl_negate_bit_ati = int(0x00000004)
	gl_bias_bit_ati   = int(0x00000008)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="TraceMaskMESA" type="bitmask" |>
pub const (
	gl_trace_operations_bit_mesa = int(0x0001)
	gl_trace_primitives_bit_mesa = int(0x0002)
	gl_trace_arrays_bit_mesa     = int(0x0004)
	gl_trace_textures_bit_mesa   = int(0x0008)
	gl_trace_pixels_bit_mesa     = int(0x0010)
	gl_trace_errors_bit_mesa     = int(0x0020)
	gl_trace_all_bits_mesa       = int(0xFFFF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="PathFontStyle" type="bitmask" |>
pub const (
	gl_bold_bit_nv   = int(0x01)
	gl_italic_bit_nv = int(0x02)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="PathMetricMask" type="bitmask" |>
pub const (
	gl_glyph_width_bit_nv                      = int(0x01)
	gl_glyph_height_bit_nv                     = int(0x02)
	gl_glyph_horizontal_bearing_x_bit_nv       = int(0x04)
	gl_glyph_horizontal_bearing_y_bit_nv       = int(0x08)
	gl_glyph_horizontal_bearing_advance_bit_nv = int(0x10)
	gl_glyph_vertical_bearing_x_bit_nv         = int(0x20)
	gl_glyph_vertical_bearing_y_bit_nv         = int(0x40)
	gl_glyph_vertical_bearing_advance_bit_nv   = int(0x80)
	gl_glyph_has_kerning_bit_nv                = int(0x100)
	gl_font_x_min_bounds_bit_nv                = int(0x00010000)
	gl_font_y_min_bounds_bit_nv                = int(0x00020000)
	gl_font_x_max_bounds_bit_nv                = int(0x00040000)
	gl_font_y_max_bounds_bit_nv                = int(0x00080000)
	gl_font_units_per_em_bit_nv                = int(0x00100000)
	gl_font_ascender_bit_nv                    = int(0x00200000)
	gl_font_descender_bit_nv                   = int(0x00400000)
	gl_font_height_bit_nv                      = int(0x00800000)
	gl_font_max_advance_width_bit_nv           = int(0x01000000)
	gl_font_max_advance_height_bit_nv          = int(0x02000000)
	gl_font_underline_position_bit_nv          = int(0x04000000)
	gl_font_underline_thickness_bit_nv         = int(0x08000000)
	gl_font_has_kerning_bit_nv                 = int(0x10000000)
	gl_font_num_glyph_indices_bit_nv           = int(0x20000000)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="PerformanceQueryCapsMaskINTEL" type="bitmask" |>
pub const (
	gl_perfquery_single_context_intel = int(0x00000000)
	gl_perfquery_global_context_intel = int(0x00000001)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="VertexHintsMaskPGI" type="bitmask" |>
pub const (
	gl_vertex23_bit_pgi                = int(0x00000004)
	gl_vertex4_bit_pgi                 = int(0x00000008)
	gl_color3_bit_pgi                  = int(0x00010000)
	gl_color4_bit_pgi                  = int(0x00020000)
	gl_edgeflag_bit_pgi                = int(0x00040000)
	gl_index_bit_pgi                   = int(0x00080000)
	gl_mat_ambient_bit_pgi             = int(0x00100000)
	gl_mat_ambient_and_diffuse_bit_pgi = int(0x00200000)
	gl_mat_diffuse_bit_pgi             = int(0x00400000)
	gl_mat_emission_bit_pgi            = int(0x00800000)
	gl_mat_color_indexes_bit_pgi       = int(0x01000000)
	gl_mat_shininess_bit_pgi           = int(0x02000000)
	gl_mat_specular_bit_pgi            = int(0x04000000)
	gl_normal_bit_pgi                  = int(0x08000000)
	gl_texcoord1_bit_pgi               = int(0x10000000)
	gl_texcoord2_bit_pgi               = int(0x20000000)
	gl_texcoord3_bit_pgi               = int(0x40000000)
	gl_texcoord4_bit_pgi               = int(0x80000000)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="BufferBitQCOM" type="bitmask" |>
pub const (
	gl_color_buffer_bit0_qcom       = int(0x00000001)
	gl_color_buffer_bit1_qcom       = int(0x00000002)
	gl_color_buffer_bit2_qcom       = int(0x00000004)
	gl_color_buffer_bit3_qcom       = int(0x00000008)
	gl_color_buffer_bit4_qcom       = int(0x00000010)
	gl_color_buffer_bit5_qcom       = int(0x00000020)
	gl_color_buffer_bit6_qcom       = int(0x00000040)
	gl_color_buffer_bit7_qcom       = int(0x00000080)
	gl_depth_buffer_bit0_qcom       = int(0x00000100)
	gl_depth_buffer_bit1_qcom       = int(0x00000200)
	gl_depth_buffer_bit2_qcom       = int(0x00000400)
	gl_depth_buffer_bit3_qcom       = int(0x00000800)
	gl_depth_buffer_bit4_qcom       = int(0x00001000)
	gl_depth_buffer_bit5_qcom       = int(0x00002000)
	gl_depth_buffer_bit6_qcom       = int(0x00004000)
	gl_depth_buffer_bit7_qcom       = int(0x00008000)
	gl_stencil_buffer_bit0_qcom     = int(0x00010000)
	gl_stencil_buffer_bit1_qcom     = int(0x00020000)
	gl_stencil_buffer_bit2_qcom     = int(0x00040000)
	gl_stencil_buffer_bit3_qcom     = int(0x00080000)
	gl_stencil_buffer_bit4_qcom     = int(0x00100000)
	gl_stencil_buffer_bit5_qcom     = int(0x00200000)
	gl_stencil_buffer_bit6_qcom     = int(0x00400000)
	gl_stencil_buffer_bit7_qcom     = int(0x00800000)
	gl_multisample_buffer_bit0_qcom = int(0x01000000)
	gl_multisample_buffer_bit1_qcom = int(0x02000000)
	gl_multisample_buffer_bit2_qcom = int(0x04000000)
	gl_multisample_buffer_bit3_qcom = int(0x08000000)
	gl_multisample_buffer_bit4_qcom = int(0x10000000)
	gl_multisample_buffer_bit5_qcom = int(0x20000000)
	gl_multisample_buffer_bit6_qcom = int(0x40000000)
	gl_multisample_buffer_bit7_qcom = int(0x80000000)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="FoveationConfigBitQCOM" type="bitmask" |>
pub const (
	gl_foveation_enable_bit_qcom                   = int(0x00000001)
	gl_foveation_scaled_bin_method_bit_qcom        = int(0x00000002)
	gl_foveation_subsampled_layout_method_bit_qcom = int(0x00000004)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="FfdMaskSGIX" type="bitmask" |>
pub const (
	gl_texture_deformation_bit_sgix  = int(0x00000001)
	gl_geometry_deformation_bit_sgix = int(0x00000002)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="CommandOpcodesNV" vendor="NV" comment="For NV_command_list." |>
pub const (
	gl_terminate_sequence_command_nv      = int(0x0000)
	gl_nop_command_nv                     = int(0x0001)
	gl_draw_elements_command_nv           = int(0x0002)
	gl_draw_arrays_command_nv             = int(0x0003)
	gl_draw_elements_strip_command_nv     = int(0x0004)
	gl_draw_arrays_strip_command_nv       = int(0x0005)
	gl_draw_elements_instanced_command_nv = int(0x0006)
	gl_draw_arrays_instanced_command_nv   = int(0x0007)
	gl_element_address_command_nv         = int(0x0008)
	gl_attribute_address_command_nv       = int(0x0009)
	gl_uniform_address_command_nv         = int(0x000A)
	gl_blend_color_command_nv             = int(0x000B)
	gl_stencil_ref_command_nv             = int(0x000C)
	gl_line_width_command_nv              = int(0x000D)
	gl_polygon_offset_command_nv          = int(0x000E)
	gl_alpha_ref_command_nv               = int(0x000F)
	gl_viewport_command_nv                = int(0x0010)
	gl_scissor_command_nv                 = int(0x0011)
	gl_front_face_command_nv              = int(0x0012)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="MapTextureFormatINTEL" vendor="INTEL" comment="Texture memory layouts for INTEL_map_texture" |>
pub const (
	gl_layout_default_intel           = int(0)
	gl_layout_linear_intel            = int(1)
	gl_layout_linear_cpu_cached_intel = int(2)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="PathRenderingTokenNV" vendor="NV" |>
pub const (
	gl_close_path_nv                         = int(0x00)
	gl_move_to_nv                            = int(0x02)
	gl_relative_move_to_nv                   = int(0x03)
	gl_line_to_nv                            = int(0x04)
	gl_relative_line_to_nv                   = int(0x05)
	gl_horizontal_line_to_nv                 = int(0x06)
	gl_relative_horizontal_line_to_nv        = int(0x07)
	gl_vertical_line_to_nv                   = int(0x08)
	gl_relative_vertical_line_to_nv          = int(0x09)
	gl_quadratic_curve_to_nv                 = int(0x0A)
	gl_relative_quadratic_curve_to_nv        = int(0x0B)
	gl_cubic_curve_to_nv                     = int(0x0C)
	gl_relative_cubic_curve_to_nv            = int(0x0D)
	gl_smooth_quadratic_curve_to_nv          = int(0x0E)
	gl_relative_smooth_quadratic_curve_to_nv = int(0x0F)
	gl_smooth_cubic_curve_to_nv              = int(0x10)
	gl_relative_smooth_cubic_curve_to_nv     = int(0x11)
	gl_small_ccw_arc_to_nv                   = int(0x12)
	gl_relative_small_ccw_arc_to_nv          = int(0x13)
	gl_small_cw_arc_to_nv                    = int(0x14)
	gl_relative_small_cw_arc_to_nv           = int(0x15)
	gl_large_ccw_arc_to_nv                   = int(0x16)
	gl_relative_large_ccw_arc_to_nv          = int(0x17)
	gl_large_cw_arc_to_nv                    = int(0x18)
	gl_relative_large_cw_arc_to_nv           = int(0x19)
	gl_conic_curve_to_nv                     = int(0x1A)
	gl_relative_conic_curve_to_nv            = int(0x1B)
	gl_shared_edge_nv                        = int(0xC0)
	gl_rounded_rect_nv                       = int(0xE8)
	gl_relative_rounded_rect_nv              = int(0xE9)
	gl_rounded_rect2_nv                      = int(0xEA)
	gl_relative_rounded_rect2_nv             = int(0xEB)
	gl_rounded_rect4_nv                      = int(0xEC)
	gl_relative_rounded_rect4_nv             = int(0xED)
	gl_rounded_rect8_nv                      = int(0xEE)
	gl_relative_rounded_rect8_nv             = int(0xEF)
	gl_restart_path_nv                       = int(0xF0)
	gl_dup_first_cubic_curve_to_nv           = int(0xF2)
	gl_dup_last_cubic_curve_to_nv            = int(0xF4)
	gl_rect_nv                               = int(0xF6)
	gl_relative_rect_nv                      = int(0xF7)
	gl_circular_ccw_arc_to_nv                = int(0xF8)
	gl_circular_cw_arc_to_nv                 = int(0xFA)
	gl_circular_tangent_arc_to_nv            = int(0xFC)
	gl_arc_to_nv                             = int(0xFE)
	gl_relative_arc_to_nv                    = int(0xFF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="TransformFeedbackTokenNV" vendor="NV" comment="For NV_transform_feedback. No clue why small negative values are used" |>
pub const (
	gl_next_buffer_nv      = int(-2)
	gl_skip_components4_nv = int(-3)
	gl_skip_components3_nv = int(-4)
	gl_skip_components2_nv = int(-5)
	gl_skip_components1_nv = int(-6)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="TriangleListSUN" vendor="SUN" |>
pub const (
	gl_restart_sun        = int(0x0001)
	gl_replace_middle_sun = int(0x0002)
	gl_replace_oldest_sun = int(0x0003)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" group="SpecialNumbers" vendor="ARB" comment="Tokens whose numeric value is intrinsically meaningful" |>
pub const (
	gl_false                 = int(0)
	gl_no_error              = int(0)
	gl_zero                  = int(0)
	gl_none                  = int(0)
	gl_none_oes              = int(0)
	gl_true                  = int(1)
	gl_one                   = int(1)
	gl_invalid_index         = int(0xFFFFFFFF)
	gl_all_pixels_amd        = int(0xFFFFFFFF)
	gl_timeout_ignored       = int(0xFFFFFFFFFFFFFFFF)
	gl_timeout_ignored_apple = int(0xFFFFFFFFFFFFFFFF)
	gl_version_es_cl_1_0     = int(1)
	gl_version_es_cm_1_1     = int(1)
	gl_version_es_cl_1_1     = int(1)
	gl_uuid_size_ext         = int(16)
	gl_luid_size_ext         = int(8)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x0000" end="0x7FFF" vendor="ARB" comment="Mostly OpenGL 1.0/1.1 enum assignments. Unused ranges should generally remain unused." |>
pub const (
	gl_points                             = int(0x0000)
	gl_lines                              = int(0x0001)
	gl_line_loop                          = int(0x0002)
	gl_line_strip                         = int(0x0003)
	gl_triangles                          = int(0x0004)
	gl_triangle_strip                     = int(0x0005)
	gl_triangle_fan                       = int(0x0006)
	gl_quads                              = int(0x0007)
	gl_quads_ext                          = int(0x0007)
	gl_quads_oes                          = int(0x0007)
	gl_quad_strip                         = int(0x0008)
	gl_polygon                            = int(0x0009)
	gl_lines_adjacency                    = int(0x000A)
	gl_lines_adjacency_arb                = int(0x000A)
	gl_lines_adjacency_ext                = int(0x000A)
	gl_lines_adjacency_oes                = int(0x000A)
	gl_line_strip_adjacency               = int(0x000B)
	gl_line_strip_adjacency_arb           = int(0x000B)
	gl_line_strip_adjacency_ext           = int(0x000B)
	gl_line_strip_adjacency_oes           = int(0x000B)
	gl_triangles_adjacency                = int(0x000C)
	gl_triangles_adjacency_arb            = int(0x000C)
	gl_triangles_adjacency_ext            = int(0x000C)
	gl_triangles_adjacency_oes            = int(0x000C)
	gl_triangle_strip_adjacency           = int(0x000D)
	gl_triangle_strip_adjacency_arb       = int(0x000D)
	gl_triangle_strip_adjacency_ext       = int(0x000D)
	gl_triangle_strip_adjacency_oes       = int(0x000D)
	gl_patches                            = int(0x000E)
	gl_patches_ext                        = int(0x000E)
	gl_patches_oes                        = int(0x000E)
	gl_accum                              = int(0x0100)
	gl_load                               = int(0x0101)
	gl_return                             = int(0x0102)
	gl_mult                               = int(0x0103)
	gl_add                                = int(0x0104)
	gl_never                              = int(0x0200)
	gl_less                               = int(0x0201)
	gl_equal                              = int(0x0202)
	gl_lequal                             = int(0x0203)
	gl_greater                            = int(0x0204)
	gl_notequal                           = int(0x0205)
	gl_gequal                             = int(0x0206)
	gl_always                             = int(0x0207)
	gl_src_color                          = int(0x0300)
	gl_one_minus_src_color                = int(0x0301)
	gl_src_alpha                          = int(0x0302)
	gl_one_minus_src_alpha                = int(0x0303)
	gl_dst_alpha                          = int(0x0304)
	gl_one_minus_dst_alpha                = int(0x0305)
	gl_dst_color                          = int(0x0306)
	gl_one_minus_dst_color                = int(0x0307)
	gl_src_alpha_saturate                 = int(0x0308)
	gl_src_alpha_saturate_ext             = int(0x0308)
	gl_front_left                         = int(0x0400)
	gl_front_right                        = int(0x0401)
	gl_back_left                          = int(0x0402)
	gl_back_right                         = int(0x0403)
	gl_front                              = int(0x0404)
	gl_back                               = int(0x0405)
	gl_left                               = int(0x0406)
	gl_right                              = int(0x0407)
	gl_front_and_back                     = int(0x0408)
	gl_aux0                               = int(0x0409)
	gl_aux1                               = int(0x040A)
	gl_aux2                               = int(0x040B)
	gl_aux3                               = int(0x040C)
	gl_invalid_enum                       = int(0x0500)
	gl_invalid_value                      = int(0x0501)
	gl_invalid_operation                  = int(0x0502)
	gl_stack_overflow                     = int(0x0503)
	gl_stack_overflow_khr                 = int(0x0503)
	gl_stack_underflow                    = int(0x0504)
	gl_stack_underflow_khr                = int(0x0504)
	gl_out_of_memory                      = int(0x0505)
	gl_invalid_framebuffer_operation      = int(0x0506)
	gl_invalid_framebuffer_operation_ext  = int(0x0506)
	gl_invalid_framebuffer_operation_oes  = int(0x0506)
	gl_context_lost                       = int(0x0507)
	gl_context_lost_khr                   = int(0x0507)
	gl_2d                                 = int(0x0600)
	gl_3d                                 = int(0x0601)
	gl_3d_color                           = int(0x0602)
	gl_3d_color_texture                   = int(0x0603)
	gl_4d_color_texture                   = int(0x0604)
	gl_pass_through_token                 = int(0x0700)
	gl_point_token                        = int(0x0701)
	gl_line_token                         = int(0x0702)
	gl_polygon_token                      = int(0x0703)
	gl_bitmap_token                       = int(0x0704)
	gl_draw_pixel_token                   = int(0x0705)
	gl_copy_pixel_token                   = int(0x0706)
	gl_line_reset_token                   = int(0x0707)
	gl_exp                                = int(0x0800)
	gl_exp2                               = int(0x0801)
	gl_cw                                 = int(0x0900)
	gl_ccw                                = int(0x0901)
	gl_coeff                              = int(0x0A00)
	gl_order                              = int(0x0A01)
	gl_domain                             = int(0x0A02)
	gl_current_color                      = int(0x0B00)
	gl_current_index                      = int(0x0B01)
	gl_current_normal                     = int(0x0B02)
	gl_current_texture_coords             = int(0x0B03)
	gl_current_raster_color               = int(0x0B04)
	gl_current_raster_index               = int(0x0B05)
	gl_current_raster_texture_coords      = int(0x0B06)
	gl_current_raster_position            = int(0x0B07)
	gl_current_raster_position_valid      = int(0x0B08)
	gl_current_raster_distance            = int(0x0B09)
	gl_point_smooth                       = int(0x0B10)
	gl_point_size                         = int(0x0B11)
	gl_point_size_range                   = int(0x0B12)
	gl_smooth_point_size_range            = int(0x0B12)
	gl_point_size_granularity             = int(0x0B13)
	gl_smooth_point_size_granularity      = int(0x0B13)
	gl_line_smooth                        = int(0x0B20)
	gl_line_width                         = int(0x0B21)
	gl_line_width_range                   = int(0x0B22)
	gl_smooth_line_width_range            = int(0x0B22)
	gl_line_width_granularity             = int(0x0B23)
	gl_smooth_line_width_granularity      = int(0x0B23)
	gl_line_stipple                       = int(0x0B24)
	gl_line_stipple_pattern               = int(0x0B25)
	gl_line_stipple_repeat                = int(0x0B26)
	gl_list_mode                          = int(0x0B30)
	gl_max_list_nesting                   = int(0x0B31)
	gl_list_base                          = int(0x0B32)
	gl_list_index                         = int(0x0B33)
	gl_polygon_mode                       = int(0x0B40)
	gl_polygon_mode_nv                    = int(0x0B40)
	gl_polygon_smooth                     = int(0x0B41)
	gl_polygon_stipple                    = int(0x0B42)
	gl_edge_flag                          = int(0x0B43)
	gl_cull_face_const                    = int(0x0B44) // because its also a function
	gl_cull_face_mode                     = int(0x0B45)
	gl_front_face                         = int(0x0B46)
	gl_lighting                           = int(0x0B50)
	gl_light_model_local_viewer           = int(0x0B51)
	gl_light_model_two_side               = int(0x0B52)
	gl_light_model_ambient                = int(0x0B53)
	gl_shade_model                        = int(0x0B54)
	gl_color_material_face                = int(0x0B55)
	gl_color_material_parameter           = int(0x0B56)
	gl_color_material                     = int(0x0B57)
	gl_fog                                = int(0x0B60)
	gl_fog_index                          = int(0x0B61)
	gl_fog_density                        = int(0x0B62)
	gl_fog_start                          = int(0x0B63)
	gl_fog_end                            = int(0x0B64)
	gl_fog_mode                           = int(0x0B65)
	gl_fog_color                          = int(0x0B66)
	gl_depth_range                        = int(0x0B70)
	gl_depth_test                         = int(0x0B71)
	gl_depth_writemask                    = int(0x0B72)
	gl_depth_clear_value                  = int(0x0B73)
	gl_depth_func                         = int(0x0B74)
	gl_accum_clear_value                  = int(0x0B80)
	gl_stencil_test                       = int(0x0B90)
	gl_stencil_clear_value                = int(0x0B91)
	gl_stencil_func                       = int(0x0B92)
	gl_stencil_value_mask                 = int(0x0B93)
	gl_stencil_fail                       = int(0x0B94)
	gl_stencil_pass_depth_fail            = int(0x0B95)
	gl_stencil_pass_depth_pass            = int(0x0B96)
	gl_stencil_ref                        = int(0x0B97)
	gl_stencil_writemask                  = int(0x0B98)
	gl_matrix_mode                        = int(0x0BA0)
	gl_normalize                          = int(0x0BA1)
	gl_viewport                           = int(0x0BA2)
	gl_modelview_stack_depth              = int(0x0BA3)
	gl_modelview0_stack_depth_ext         = int(0x0BA3)
	gl_path_modelview_stack_depth_nv      = int(0x0BA3)
	gl_projection_stack_depth             = int(0x0BA4)
	gl_path_projection_stack_depth_nv     = int(0x0BA4)
	gl_texture_stack_depth                = int(0x0BA5)
	gl_modelview_matrix                   = int(0x0BA6)
	gl_modelview0_matrix_ext              = int(0x0BA6)
	gl_path_modelview_matrix_nv           = int(0x0BA6)
	gl_projection_matrix                  = int(0x0BA7)
	gl_path_projection_matrix_nv          = int(0x0BA7)
	gl_texture_matrix                     = int(0x0BA8)
	gl_attrib_stack_depth                 = int(0x0BB0)
	gl_client_attrib_stack_depth          = int(0x0BB1)
	gl_alpha_test                         = int(0x0BC0)
	gl_alpha_test_qcom                    = int(0x0BC0)
	gl_alpha_test_func                    = int(0x0BC1)
	gl_alpha_test_func_qcom               = int(0x0BC1)
	gl_alpha_test_ref                     = int(0x0BC2)
	gl_alpha_test_ref_qcom                = int(0x0BC2)
	gl_dither                             = int(0x0BD0)
	gl_blend_dst                          = int(0x0BE0)
	gl_blend_src                          = int(0x0BE1)
	gl_blend                              = int(0x0BE2)
	gl_logic_op_mode                      = int(0x0BF0)
	gl_index_logic_op                     = int(0x0BF1)
	gl_logic_op                           = int(0x0BF1)
	gl_color_logic_op                     = int(0x0BF2)
	gl_aux_buffers                        = int(0x0C00)
	gl_draw_buffer                        = int(0x0C01)
	gl_draw_buffer_ext                    = int(0x0C01)
	gl_read_buffer                        = int(0x0C02)
	gl_read_buffer_ext                    = int(0x0C02)
	gl_read_buffer_nv                     = int(0x0C02)
	gl_scissor_box                        = int(0x0C10)
	gl_scissor_test                       = int(0x0C11)
	gl_index_clear_value                  = int(0x0C20)
	gl_index_writemask                    = int(0x0C21)
	gl_color_clear_value                  = int(0x0C22)
	gl_color_writemask                    = int(0x0C23)
	gl_index_mode                         = int(0x0C30)
	gl_rgba_mode                          = int(0x0C31)
	gl_doublebuffer                       = int(0x0C32)
	gl_stereo                             = int(0x0C33)
	gl_render_mode                        = int(0x0C40)
	gl_perspective_correction_hint        = int(0x0C50)
	gl_point_smooth_hint                  = int(0x0C51)
	gl_line_smooth_hint                   = int(0x0C52)
	gl_polygon_smooth_hint                = int(0x0C53)
	gl_fog_hint                           = int(0x0C54)
	gl_texture_gen_s                      = int(0x0C60)
	gl_texture_gen_t                      = int(0x0C61)
	gl_texture_gen_r                      = int(0x0C62)
	gl_texture_gen_q                      = int(0x0C63)
	gl_pixel_map_i_to_i                   = int(0x0C70)
	gl_pixel_map_s_to_s                   = int(0x0C71)
	gl_pixel_map_i_to_r                   = int(0x0C72)
	gl_pixel_map_i_to_g                   = int(0x0C73)
	gl_pixel_map_i_to_b                   = int(0x0C74)
	gl_pixel_map_i_to_a                   = int(0x0C75)
	gl_pixel_map_r_to_r                   = int(0x0C76)
	gl_pixel_map_g_to_g                   = int(0x0C77)
	gl_pixel_map_b_to_b                   = int(0x0C78)
	gl_pixel_map_a_to_a                   = int(0x0C79)
	gl_pixel_map_i_to_i_size              = int(0x0CB0)
	gl_pixel_map_s_to_s_size              = int(0x0CB1)
	gl_pixel_map_i_to_r_size              = int(0x0CB2)
	gl_pixel_map_i_to_g_size              = int(0x0CB3)
	gl_pixel_map_i_to_b_size              = int(0x0CB4)
	gl_pixel_map_i_to_a_size              = int(0x0CB5)
	gl_pixel_map_r_to_r_size              = int(0x0CB6)
	gl_pixel_map_g_to_g_size              = int(0x0CB7)
	gl_pixel_map_b_to_b_size              = int(0x0CB8)
	gl_pixel_map_a_to_a_size              = int(0x0CB9)
	gl_unpack_swap_bytes                  = int(0x0CF0)
	gl_unpack_lsb_first                   = int(0x0CF1)
	gl_unpack_row_length                  = int(0x0CF2)
	gl_unpack_row_length_ext              = int(0x0CF2)
	gl_unpack_skip_rows                   = int(0x0CF3)
	gl_unpack_skip_rows_ext               = int(0x0CF3)
	gl_unpack_skip_pixels                 = int(0x0CF4)
	gl_unpack_skip_pixels_ext             = int(0x0CF4)
	gl_unpack_alignment                   = int(0x0CF5)
	gl_pack_swap_bytes                    = int(0x0D00)
	gl_pack_lsb_first                     = int(0x0D01)
	gl_pack_row_length                    = int(0x0D02)
	gl_pack_row_length_nv                 = int(0x0D02)
	gl_pack_skip_rows                     = int(0x0D03)
	gl_pack_skip_rows_nv                  = int(0x0D03)
	gl_pack_skip_pixels                   = int(0x0D04)
	gl_pack_skip_pixels_nv                = int(0x0D04)
	gl_pack_alignment                     = int(0x0D05)
	gl_map_color                          = int(0x0D10)
	gl_map_stencil                        = int(0x0D11)
	gl_index_shift                        = int(0x0D12)
	gl_index_offset                       = int(0x0D13)
	gl_red_scale                          = int(0x0D14)
	gl_red_bias                           = int(0x0D15)
	gl_zoom_x                             = int(0x0D16)
	gl_zoom_y                             = int(0x0D17)
	gl_green_scale                        = int(0x0D18)
	gl_green_bias                         = int(0x0D19)
	gl_blue_scale                         = int(0x0D1A)
	gl_blue_bias                          = int(0x0D1B)
	gl_alpha_scale                        = int(0x0D1C)
	gl_alpha_bias                         = int(0x0D1D)
	gl_depth_scale                        = int(0x0D1E)
	gl_depth_bias                         = int(0x0D1F)
	gl_max_eval_order                     = int(0x0D30)
	gl_max_lights                         = int(0x0D31)
	gl_max_clip_planes                    = int(0x0D32)
	gl_max_clip_planes_img                = int(0x0D32)
	gl_max_clip_distances                 = int(0x0D32)
	gl_max_clip_distances_ext             = int(0x0D32)
	gl_max_clip_distances_apple           = int(0x0D32)
	gl_max_texture_size                   = int(0x0D33)
	gl_max_pixel_map_table                = int(0x0D34)
	gl_max_attrib_stack_depth             = int(0x0D35)
	gl_max_modelview_stack_depth          = int(0x0D36)
	gl_path_max_modelview_stack_depth_nv  = int(0x0D36)
	gl_max_name_stack_depth               = int(0x0D37)
	gl_max_projection_stack_depth         = int(0x0D38)
	gl_path_max_projection_stack_depth_nv = int(0x0D38)
	gl_max_texture_stack_depth            = int(0x0D39)
	gl_max_viewport_dims                  = int(0x0D3A)
	gl_max_client_attrib_stack_depth      = int(0x0D3B)
	gl_subpixel_bits                      = int(0x0D50)
	gl_index_bits                         = int(0x0D51)
	gl_red_bits                           = int(0x0D52)
	gl_green_bits                         = int(0x0D53)
	gl_blue_bits                          = int(0x0D54)
	gl_alpha_bits                         = int(0x0D55)
	gl_depth_bits                         = int(0x0D56)
	gl_stencil_bits                       = int(0x0D57)
	gl_accum_red_bits                     = int(0x0D58)
	gl_accum_green_bits                   = int(0x0D59)
	gl_accum_blue_bits                    = int(0x0D5A)
	gl_accum_alpha_bits                   = int(0x0D5B)
	gl_name_stack_depth                   = int(0x0D70)
	gl_auto_normal                        = int(0x0D80)
	gl_map1_color_4                       = int(0x0D90)
	gl_map1_index                         = int(0x0D91)
	gl_map1_normal                        = int(0x0D92)
	gl_map1_texture_coord_1               = int(0x0D93)
	gl_map1_texture_coord_2               = int(0x0D94)
	gl_map1_texture_coord_3               = int(0x0D95)
	gl_map1_texture_coord_4               = int(0x0D96)
	gl_map1_vertex_3                      = int(0x0D97)
	gl_map1_vertex_4                      = int(0x0D98)
	gl_map2_color_4                       = int(0x0DB0)
	gl_map2_index                         = int(0x0DB1)
	gl_map2_normal                        = int(0x0DB2)
	gl_map2_texture_coord_1               = int(0x0DB3)
	gl_map2_texture_coord_2               = int(0x0DB4)
	gl_map2_texture_coord_3               = int(0x0DB5)
	gl_map2_texture_coord_4               = int(0x0DB6)
	gl_map2_vertex_3                      = int(0x0DB7)
	gl_map2_vertex_4                      = int(0x0DB8)
	gl_map1_grid_domain                   = int(0x0DD0)
	gl_map1_grid_segments                 = int(0x0DD1)
	gl_map2_grid_domain                   = int(0x0DD2)
	gl_map2_grid_segments                 = int(0x0DD3)
	gl_texture_1d                         = int(0x0DE0)
	gl_texture_2d                         = int(0x0DE1)
	gl_feedback_buffer_pointer            = int(0x0DF0)
	gl_feedback_buffer_size               = int(0x0DF1)
	gl_feedback_buffer_type               = int(0x0DF2)
	gl_selection_buffer_pointer           = int(0x0DF3)
	gl_selection_buffer_size              = int(0x0DF4)
	gl_texture_width                      = int(0x1000)
	gl_texture_height                     = int(0x1001)
	gl_texture_internal_format            = int(0x1003)
	gl_texture_components                 = int(0x1003)
	gl_texture_border_color               = int(0x1004)
	gl_texture_border_color_ext           = int(0x1004)
	gl_texture_border_color_nv            = int(0x1004)
	gl_texture_border_color_oes           = int(0x1004)
	gl_texture_border                     = int(0x1005)
	gl_texture_target                     = int(0x1006)
	gl_dont_care                          = int(0x1100)
	gl_fastest                            = int(0x1101)
	gl_nicest                             = int(0x1102)
	gl_ambient                            = int(0x1200)
	gl_diffuse                            = int(0x1201)
	gl_specular                           = int(0x1202)
	gl_position                           = int(0x1203)
	gl_spot_direction                     = int(0x1204)
	gl_spot_exponent                      = int(0x1205)
	gl_spot_cutoff                        = int(0x1206)
	gl_constant_attenuation               = int(0x1207)
	gl_linear_attenuation                 = int(0x1208)
	gl_quadratic_attenuation              = int(0x1209)
	gl_compile                            = int(0x1300)
	gl_compile_and_execute                = int(0x1301)
	gl_byte                               = int(0x1400)
	gl_unsigned_byte                      = int(0x1401)
	gl_short                              = int(0x1402)
	gl_unsigned_short                     = int(0x1403)
	gl_int                                = int(0x1404)
	gl_unsigned_int                       = int(0x1405)
	gl_float                              = int(0x1406)
	gl_2_bytes                            = int(0x1407)
	gl_2_bytes_nv                         = int(0x1407)
	gl_3_bytes                            = int(0x1408)
	gl_3_bytes_nv                         = int(0x1408)
	gl_4_bytes                            = int(0x1409)
	gl_4_bytes_nv                         = int(0x1409)
	gl_double                             = int(0x140A)
	gl_double_ext                         = int(0x140A)
	gl_half_float                         = int(0x140B)
	gl_half_float_arb                     = int(0x140B)
	gl_half_float_nv                      = int(0x140B)
	gl_half_apple                         = int(0x140B)
	gl_fixed                              = int(0x140C)
	gl_fixed_oes                          = int(0x140C)
	gl_int64_arb                          = int(0x140E)
	gl_int64_nv                           = int(0x140E)
	gl_unsigned_int64_arb                 = int(0x140F)
	gl_unsigned_int64_nv                  = int(0x140F)
	gl_clear                              = int(0x1500)
	gl_and                                = int(0x1501)
	gl_and_reverse                        = int(0x1502)
	gl_copy                               = int(0x1503)
	gl_and_inverted                       = int(0x1504)
	gl_noop                               = int(0x1505)
	gl_xor                                = int(0x1506)
	gl_xor_nv                             = int(0x1506)
	gl_or                                 = int(0x1507)
	gl_nor                                = int(0x1508)
	gl_equiv                              = int(0x1509)
	gl_invert                             = int(0x150A)
	gl_or_reverse                         = int(0x150B)
	gl_copy_inverted                      = int(0x150C)
	gl_or_inverted                        = int(0x150D)
	gl_nand                               = int(0x150E)
	gl_set                                = int(0x150F)
	gl_emission                           = int(0x1600)
	gl_shininess                          = int(0x1601)
	gl_ambient_and_diffuse                = int(0x1602)
	gl_color_indexes                      = int(0x1603)
	gl_modelview                          = int(0x1700)
	gl_modelview0_arb                     = int(0x1700)
	gl_modelview0_ext                     = int(0x1700)
	gl_path_modelview_nv                  = int(0x1700)
	gl_projection                         = int(0x1701)
	gl_path_projection_nv                 = int(0x1701)
	gl_texture                            = int(0x1702)
	gl_color                              = int(0x1800)
	gl_color_ext                          = int(0x1800)
	gl_depth                              = int(0x1801)
	gl_depth_ext                          = int(0x1801)
	gl_stencil                            = int(0x1802)
	gl_stencil_ext                        = int(0x1802)
	gl_color_index                        = int(0x1900)
	gl_stencil_index                      = int(0x1901)
	gl_stencil_index_oes                  = int(0x1901)
	gl_depth_component                    = int(0x1902)
	gl_red                                = int(0x1903)
	gl_red_ext                            = int(0x1903)
	gl_red_nv                             = int(0x1903)
	gl_green                              = int(0x1904)
	gl_green_nv                           = int(0x1904)
	gl_blue                               = int(0x1905)
	gl_blue_nv                            = int(0x1905)
	gl_alpha                              = int(0x1906)
	gl_rgb                                = int(0x1907)
	gl_rgba                               = int(0x1908)
	gl_luminance                          = int(0x1909)
	gl_luminance_alpha                    = int(0x190A)
	gl_bitmap                             = int(0x1A00)
	gl_point                              = int(0x1B00)
	gl_point_nv                           = int(0x1B00)
	gl_line                               = int(0x1B01)
	gl_line_nv                            = int(0x1B01)
	gl_fill                               = int(0x1B02)
	gl_fill_nv                            = int(0x1B02)
	gl_render                             = int(0x1C00)
	gl_feedback                           = int(0x1C01)
	gl_select                             = int(0x1C02)
	gl_flat                               = int(0x1D00)
	gl_smooth                             = int(0x1D01)
	gl_keep                               = int(0x1E00)
	gl_replace                            = int(0x1E01)
	gl_incr                               = int(0x1E02)
	gl_decr                               = int(0x1E03)
	gl_vendor                             = int(0x1F00)
	gl_renderer                           = int(0x1F01)
	gl_version                            = int(0x1F02)
	gl_extensions                         = int(0x1F03)
	gl_s                                  = int(0x2000)
	gl_t                                  = int(0x2001)
	gl_r                                  = int(0x2002)
	gl_q                                  = int(0x2003)
	gl_modulate                           = int(0x2100)
	gl_decal                              = int(0x2101)
	gl_texture_env_mode                   = int(0x2200)
	gl_texture_env_color                  = int(0x2201)
	gl_texture_env                        = int(0x2300)
	gl_eye_linear                         = int(0x2400)
	gl_eye_linear_nv                      = int(0x2400)
	gl_object_linear                      = int(0x2401)
	gl_object_linear_nv                   = int(0x2401)
	gl_sphere_map                         = int(0x2402)
	gl_texture_gen_mode                   = int(0x2500)
	gl_texture_gen_mode_oes               = int(0x2500)
	gl_object_plane                       = int(0x2501)
	gl_eye_plane                          = int(0x2502)
	gl_nearest                            = int(0x2600)
	gl_linear                             = int(0x2601)
	gl_nearest_mipmap_nearest             = int(0x2700)
	gl_linear_mipmap_nearest              = int(0x2701)
	gl_nearest_mipmap_linear              = int(0x2702)
	gl_linear_mipmap_linear               = int(0x2703)
	gl_texture_mag_filter                 = int(0x2800)
	gl_texture_min_filter                 = int(0x2801)
	gl_texture_wrap_s                     = int(0x2802)
	gl_texture_wrap_t                     = int(0x2803)
	gl_clamp                              = int(0x2900)
	gl_repeat                             = int(0x2901)
	gl_polygon_offset_units               = int(0x2A00)
	gl_polygon_offset_point               = int(0x2A01)
	gl_polygon_offset_point_nv            = int(0x2A01)
	gl_polygon_offset_line                = int(0x2A02)
	gl_polygon_offset_line_nv             = int(0x2A02)
	gl_r3_g3_b2                           = int(0x2A10)
	gl_v2f                                = int(0x2A20)
	gl_v3f                                = int(0x2A21)
	gl_c4ub_v2f                           = int(0x2A22)
	gl_c4ub_v3f                           = int(0x2A23)
	gl_c3f_v3f                            = int(0x2A24)
	gl_n3f_v3f                            = int(0x2A25)
	gl_c4f_n3f_v3f                        = int(0x2A26)
	gl_t2f_v3f                            = int(0x2A27)
	gl_t4f_v4f                            = int(0x2A28)
	gl_t2f_c4ub_v3f                       = int(0x2A29)
	gl_t2f_c3f_v3f                        = int(0x2A2A)
	gl_t2f_n3f_v3f                        = int(0x2A2B)
	gl_t2f_c4f_n3f_v3f                    = int(0x2A2C)
	gl_t4f_c4f_n3f_v4f                    = int(0x2A2D)
	gl_clip_plane0                        = int(0x3000)
	gl_clip_plane0_img                    = int(0x3000)
	gl_clip_distance0                     = int(0x3000)
	gl_clip_distance0_ext                 = int(0x3000)
	gl_clip_distance0_apple               = int(0x3000)
	gl_clip_plane1                        = int(0x3001)
	gl_clip_plane1_img                    = int(0x3001)
	gl_clip_distance1                     = int(0x3001)
	gl_clip_distance1_ext                 = int(0x3001)
	gl_clip_distance1_apple               = int(0x3001)
	gl_clip_plane2                        = int(0x3002)
	gl_clip_plane2_img                    = int(0x3002)
	gl_clip_distance2                     = int(0x3002)
	gl_clip_distance2_ext                 = int(0x3002)
	gl_clip_distance2_apple               = int(0x3002)
	gl_clip_plane3                        = int(0x3003)
	gl_clip_plane3_img                    = int(0x3003)
	gl_clip_distance3                     = int(0x3003)
	gl_clip_distance3_ext                 = int(0x3003)
	gl_clip_distance3_apple               = int(0x3003)
	gl_clip_plane4                        = int(0x3004)
	gl_clip_plane4_img                    = int(0x3004)
	gl_clip_distance4                     = int(0x3004)
	gl_clip_distance4_ext                 = int(0x3004)
	gl_clip_distance4_apple               = int(0x3004)
	gl_clip_plane5                        = int(0x3005)
	gl_clip_plane5_img                    = int(0x3005)
	gl_clip_distance5                     = int(0x3005)
	gl_clip_distance5_ext                 = int(0x3005)
	gl_clip_distance5_apple               = int(0x3005)
	gl_clip_distance6                     = int(0x3006)
	gl_clip_distance6_ext                 = int(0x3006)
	gl_clip_distance6_apple               = int(0x3006)
	gl_clip_distance7                     = int(0x3007)
	gl_clip_distance7_ext                 = int(0x3007)
	gl_clip_distance7_apple               = int(0x3007)
	gl_light0                             = int(0x4000)
	gl_light1                             = int(0x4001)
	gl_light2                             = int(0x4002)
	gl_light3                             = int(0x4003)
	gl_light4                             = int(0x4004)
	gl_light5                             = int(0x4005)
	gl_light6                             = int(0x4006)
	gl_light7                             = int(0x4007)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8000" end="0x80BF" vendor="ARB" comment="The primary GL enumerant space begins here. All modern enum allocations are in this range. These enums are mostly assigned the default class since it's a great deal of not very useful work to be more specific" |>
pub const (
	gl_abgr_ext                          = int(0x8000)
	gl_constant_color                    = int(0x8001)
	gl_constant_color_ext                = int(0x8001)
	gl_one_minus_constant_color          = int(0x8002)
	gl_one_minus_constant_color_ext      = int(0x8002)
	gl_constant_alpha                    = int(0x8003)
	gl_constant_alpha_ext                = int(0x8003)
	gl_one_minus_constant_alpha          = int(0x8004)
	gl_one_minus_constant_alpha_ext      = int(0x8004)
	gl_blend_color                       = int(0x8005)
	gl_blend_color_ext                   = int(0x8005)
	gl_func_add                          = int(0x8006)
	gl_func_add_ext                      = int(0x8006)
	gl_func_add_oes                      = int(0x8006)
	gl_min                               = int(0x8007)
	gl_min_ext                           = int(0x8007)
	gl_max                               = int(0x8008)
	gl_max_ext                           = int(0x8008)
	gl_blend_equation                    = int(0x8009)
	gl_blend_equation_ext                = int(0x8009)
	gl_blend_equation_oes                = int(0x8009)
	gl_blend_equation_rgb                = int(0x8009)
	gl_blend_equation_rgb_ext            = int(0x8009)
	gl_blend_equation_rgb_oes            = int(0x8009)
	gl_func_subtract                     = int(0x800A)
	gl_func_subtract_ext                 = int(0x800A)
	gl_func_subtract_oes                 = int(0x800A)
	gl_func_reverse_subtract             = int(0x800B)
	gl_func_reverse_subtract_ext         = int(0x800B)
	gl_func_reverse_subtract_oes         = int(0x800B)
	gl_cmyk_ext                          = int(0x800C)
	gl_cmyka_ext                         = int(0x800D)
	gl_pack_cmyk_hint_ext                = int(0x800E)
	gl_unpack_cmyk_hint_ext              = int(0x800F)
	gl_convolution_1d                    = int(0x8010)
	gl_convolution_1d_ext                = int(0x8010)
	gl_convolution_2d                    = int(0x8011)
	gl_convolution_2d_ext                = int(0x8011)
	gl_separable_2d                      = int(0x8012)
	gl_separable_2d_ext                  = int(0x8012)
	gl_convolution_border_mode           = int(0x8013)
	gl_convolution_border_mode_ext       = int(0x8013)
	gl_convolution_filter_scale          = int(0x8014)
	gl_convolution_filter_scale_ext      = int(0x8014)
	gl_convolution_filter_bias           = int(0x8015)
	gl_convolution_filter_bias_ext       = int(0x8015)
	gl_reduce                            = int(0x8016)
	gl_reduce_ext                        = int(0x8016)
	gl_convolution_format                = int(0x8017)
	gl_convolution_format_ext            = int(0x8017)
	gl_convolution_width                 = int(0x8018)
	gl_convolution_width_ext             = int(0x8018)
	gl_convolution_height                = int(0x8019)
	gl_convolution_height_ext            = int(0x8019)
	gl_max_convolution_width             = int(0x801A)
	gl_max_convolution_width_ext         = int(0x801A)
	gl_max_convolution_height            = int(0x801B)
	gl_max_convolution_height_ext        = int(0x801B)
	gl_post_convolution_red_scale        = int(0x801C)
	gl_post_convolution_red_scale_ext    = int(0x801C)
	gl_post_convolution_green_scale      = int(0x801D)
	gl_post_convolution_green_scale_ext  = int(0x801D)
	gl_post_convolution_blue_scale       = int(0x801E)
	gl_post_convolution_blue_scale_ext   = int(0x801E)
	gl_post_convolution_alpha_scale      = int(0x801F)
	gl_post_convolution_alpha_scale_ext  = int(0x801F)
	gl_post_convolution_red_bias         = int(0x8020)
	gl_post_convolution_red_bias_ext     = int(0x8020)
	gl_post_convolution_green_bias       = int(0x8021)
	gl_post_convolution_green_bias_ext   = int(0x8021)
	gl_post_convolution_blue_bias        = int(0x8022)
	gl_post_convolution_blue_bias_ext    = int(0x8022)
	gl_post_convolution_alpha_bias       = int(0x8023)
	gl_post_convolution_alpha_bias_ext   = int(0x8023)
	gl_histogram                         = int(0x8024)
	gl_histogram_ext                     = int(0x8024)
	gl_proxy_histogram                   = int(0x8025)
	gl_proxy_histogram_ext               = int(0x8025)
	gl_histogram_width                   = int(0x8026)
	gl_histogram_width_ext               = int(0x8026)
	gl_histogram_format                  = int(0x8027)
	gl_histogram_format_ext              = int(0x8027)
	gl_histogram_red_size                = int(0x8028)
	gl_histogram_red_size_ext            = int(0x8028)
	gl_histogram_green_size              = int(0x8029)
	gl_histogram_green_size_ext          = int(0x8029)
	gl_histogram_blue_size               = int(0x802A)
	gl_histogram_blue_size_ext           = int(0x802A)
	gl_histogram_alpha_size              = int(0x802B)
	gl_histogram_alpha_size_ext          = int(0x802B)
	gl_histogram_luminance_size          = int(0x802C)
	gl_histogram_luminance_size_ext      = int(0x802C)
	gl_histogram_sink                    = int(0x802D)
	gl_histogram_sink_ext                = int(0x802D)
	gl_minmax                            = int(0x802E)
	gl_minmax_ext                        = int(0x802E)
	gl_minmax_format                     = int(0x802F)
	gl_minmax_format_ext                 = int(0x802F)
	gl_minmax_sink                       = int(0x8030)
	gl_minmax_sink_ext                   = int(0x8030)
	gl_table_too_large_ext               = int(0x8031)
	gl_table_too_large                   = int(0x8031)
	gl_unsigned_byte_3_3_2               = int(0x8032)
	gl_unsigned_byte_3_3_2_ext           = int(0x8032)
	gl_unsigned_short_4_4_4_4            = int(0x8033)
	gl_unsigned_short_4_4_4_4_ext        = int(0x8033)
	gl_unsigned_short_5_5_5_1            = int(0x8034)
	gl_unsigned_short_5_5_5_1_ext        = int(0x8034)
	gl_unsigned_int_8_8_8_8              = int(0x8035)
	gl_unsigned_int_8_8_8_8_ext          = int(0x8035)
	gl_unsigned_int_10_10_10_2           = int(0x8036)
	gl_unsigned_int_10_10_10_2_ext       = int(0x8036)
	gl_polygon_offset_ext                = int(0x8037)
	gl_polygon_offset_fill               = int(0x8037)
	gl_polygon_offset_factor             = int(0x8038)
	gl_polygon_offset_factor_ext         = int(0x8038)
	gl_polygon_offset_bias_ext           = int(0x8039)
	gl_rescale_normal                    = int(0x803A)
	gl_rescale_normal_ext                = int(0x803A)
	gl_alpha4                            = int(0x803B)
	gl_alpha4_ext                        = int(0x803B)
	gl_alpha8                            = int(0x803C)
	gl_alpha8_ext                        = int(0x803C)
	gl_alpha8_oes                        = int(0x803C)
	gl_alpha12                           = int(0x803D)
	gl_alpha12_ext                       = int(0x803D)
	gl_alpha16                           = int(0x803E)
	gl_alpha16_ext                       = int(0x803E)
	gl_luminance4                        = int(0x803F)
	gl_luminance4_ext                    = int(0x803F)
	gl_luminance8                        = int(0x8040)
	gl_luminance8_ext                    = int(0x8040)
	gl_luminance8_oes                    = int(0x8040)
	gl_luminance12                       = int(0x8041)
	gl_luminance12_ext                   = int(0x8041)
	gl_luminance16                       = int(0x8042)
	gl_luminance16_ext                   = int(0x8042)
	gl_luminance4_alpha4                 = int(0x8043)
	gl_luminance4_alpha4_ext             = int(0x8043)
	gl_luminance4_alpha4_oes             = int(0x8043)
	gl_luminance6_alpha2                 = int(0x8044)
	gl_luminance6_alpha2_ext             = int(0x8044)
	gl_luminance8_alpha8                 = int(0x8045)
	gl_luminance8_alpha8_ext             = int(0x8045)
	gl_luminance8_alpha8_oes             = int(0x8045)
	gl_luminance12_alpha4                = int(0x8046)
	gl_luminance12_alpha4_ext            = int(0x8046)
	gl_luminance12_alpha12               = int(0x8047)
	gl_luminance12_alpha12_ext           = int(0x8047)
	gl_luminance16_alpha16               = int(0x8048)
	gl_luminance16_alpha16_ext           = int(0x8048)
	gl_intensity                         = int(0x8049)
	gl_intensity_ext                     = int(0x8049)
	gl_intensity4                        = int(0x804A)
	gl_intensity4_ext                    = int(0x804A)
	gl_intensity8                        = int(0x804B)
	gl_intensity8_ext                    = int(0x804B)
	gl_intensity12                       = int(0x804C)
	gl_intensity12_ext                   = int(0x804C)
	gl_intensity16                       = int(0x804D)
	gl_intensity16_ext                   = int(0x804D)
	gl_rgb2_ext                          = int(0x804E)
	gl_rgb4                              = int(0x804F)
	gl_rgb4_ext                          = int(0x804F)
	gl_rgb5                              = int(0x8050)
	gl_rgb5_ext                          = int(0x8050)
	gl_rgb8                              = int(0x8051)
	gl_rgb8_ext                          = int(0x8051)
	gl_rgb8_oes                          = int(0x8051)
	gl_rgb10                             = int(0x8052)
	gl_rgb10_ext                         = int(0x8052)
	gl_rgb12                             = int(0x8053)
	gl_rgb12_ext                         = int(0x8053)
	gl_rgb16                             = int(0x8054)
	gl_rgb16_ext                         = int(0x8054)
	gl_rgba2                             = int(0x8055)
	gl_rgba2_ext                         = int(0x8055)
	gl_rgba4                             = int(0x8056)
	gl_rgba4_ext                         = int(0x8056)
	gl_rgba4_oes                         = int(0x8056)
	gl_rgb5_a1                           = int(0x8057)
	gl_rgb5_a1_ext                       = int(0x8057)
	gl_rgb5_a1_oes                       = int(0x8057)
	gl_rgba8                             = int(0x8058)
	gl_rgba8_ext                         = int(0x8058)
	gl_rgba8_oes                         = int(0x8058)
	gl_rgb10_a2                          = int(0x8059)
	gl_rgb10_a2_ext                      = int(0x8059)
	gl_rgba12                            = int(0x805A)
	gl_rgba12_ext                        = int(0x805A)
	gl_rgba16                            = int(0x805B)
	gl_rgba16_ext                        = int(0x805B)
	gl_texture_red_size                  = int(0x805C)
	gl_texture_red_size_ext              = int(0x805C)
	gl_texture_green_size                = int(0x805D)
	gl_texture_green_size_ext            = int(0x805D)
	gl_texture_blue_size                 = int(0x805E)
	gl_texture_blue_size_ext             = int(0x805E)
	gl_texture_alpha_size                = int(0x805F)
	gl_texture_alpha_size_ext            = int(0x805F)
	gl_texture_luminance_size            = int(0x8060)
	gl_texture_luminance_size_ext        = int(0x8060)
	gl_texture_intensity_size            = int(0x8061)
	gl_texture_intensity_size_ext        = int(0x8061)
	gl_replace_ext                       = int(0x8062)
	gl_proxy_texture_1d                  = int(0x8063)
	gl_proxy_texture_1d_ext              = int(0x8063)
	gl_proxy_texture_2d                  = int(0x8064)
	gl_proxy_texture_2d_ext              = int(0x8064)
	gl_texture_too_large_ext             = int(0x8065)
	gl_texture_priority                  = int(0x8066)
	gl_texture_priority_ext              = int(0x8066)
	gl_texture_resident                  = int(0x8067)
	gl_texture_resident_ext              = int(0x8067)
	gl_texture_1d_binding_ext            = int(0x8068)
	gl_texture_binding_1d                = int(0x8068)
	gl_texture_2d_binding_ext            = int(0x8069)
	gl_texture_binding_2d                = int(0x8069)
	gl_texture_3d_binding_ext            = int(0x806A)
	gl_texture_3d_binding_oes            = int(0x806A)
	gl_texture_binding_3d                = int(0x806A)
	gl_texture_binding_3d_oes            = int(0x806A)
	gl_pack_skip_images                  = int(0x806B)
	gl_pack_skip_images_ext              = int(0x806B)
	gl_pack_image_height                 = int(0x806C)
	gl_pack_image_height_ext             = int(0x806C)
	gl_unpack_skip_images                = int(0x806D)
	gl_unpack_skip_images_ext            = int(0x806D)
	gl_unpack_image_height               = int(0x806E)
	gl_unpack_image_height_ext           = int(0x806E)
	gl_texture_3d                        = int(0x806F)
	gl_texture_3d_ext                    = int(0x806F)
	gl_texture_3d_oes                    = int(0x806F)
	gl_proxy_texture_3d                  = int(0x8070)
	gl_proxy_texture_3d_ext              = int(0x8070)
	gl_texture_depth                     = int(0x8071)
	gl_texture_depth_ext                 = int(0x8071)
	gl_texture_wrap_r                    = int(0x8072)
	gl_texture_wrap_r_ext                = int(0x8072)
	gl_texture_wrap_r_oes                = int(0x8072)
	gl_max_3d_texture_size               = int(0x8073)
	gl_max_3d_texture_size_ext           = int(0x8073)
	gl_max_3d_texture_size_oes           = int(0x8073)
	gl_vertex_array                      = int(0x8074)
	gl_vertex_array_ext                  = int(0x8074)
	gl_vertex_array_khr                  = int(0x8074)
	gl_normal_array                      = int(0x8075)
	gl_normal_array_ext                  = int(0x8075)
	gl_color_array                       = int(0x8076)
	gl_color_array_ext                   = int(0x8076)
	gl_index_array                       = int(0x8077)
	gl_index_array_ext                   = int(0x8077)
	gl_texture_coord_array               = int(0x8078)
	gl_texture_coord_array_ext           = int(0x8078)
	gl_edge_flag_array                   = int(0x8079)
	gl_edge_flag_array_ext               = int(0x8079)
	gl_vertex_array_size                 = int(0x807A)
	gl_vertex_array_size_ext             = int(0x807A)
	gl_vertex_array_type                 = int(0x807B)
	gl_vertex_array_type_ext             = int(0x807B)
	gl_vertex_array_stride               = int(0x807C)
	gl_vertex_array_stride_ext           = int(0x807C)
	gl_vertex_array_count_ext            = int(0x807D)
	gl_normal_array_type                 = int(0x807E)
	gl_normal_array_type_ext             = int(0x807E)
	gl_normal_array_stride               = int(0x807F)
	gl_normal_array_stride_ext           = int(0x807F)
	gl_normal_array_count_ext            = int(0x8080)
	gl_color_array_size                  = int(0x8081)
	gl_color_array_size_ext              = int(0x8081)
	gl_color_array_type                  = int(0x8082)
	gl_color_array_type_ext              = int(0x8082)
	gl_color_array_stride                = int(0x8083)
	gl_color_array_stride_ext            = int(0x8083)
	gl_color_array_count_ext             = int(0x8084)
	gl_index_array_type                  = int(0x8085)
	gl_index_array_type_ext              = int(0x8085)
	gl_index_array_stride                = int(0x8086)
	gl_index_array_stride_ext            = int(0x8086)
	gl_index_array_count_ext             = int(0x8087)
	gl_texture_coord_array_size          = int(0x8088)
	gl_texture_coord_array_size_ext      = int(0x8088)
	gl_texture_coord_array_type          = int(0x8089)
	gl_texture_coord_array_type_ext      = int(0x8089)
	gl_texture_coord_array_stride        = int(0x808A)
	gl_texture_coord_array_stride_ext    = int(0x808A)
	gl_texture_coord_array_count_ext     = int(0x808B)
	gl_edge_flag_array_stride            = int(0x808C)
	gl_edge_flag_array_stride_ext        = int(0x808C)
	gl_edge_flag_array_count_ext         = int(0x808D)
	gl_vertex_array_pointer              = int(0x808E)
	gl_vertex_array_pointer_ext          = int(0x808E)
	gl_normal_array_pointer              = int(0x808F)
	gl_normal_array_pointer_ext          = int(0x808F)
	gl_color_array_pointer               = int(0x8090)
	gl_color_array_pointer_ext           = int(0x8090)
	gl_index_array_pointer               = int(0x8091)
	gl_index_array_pointer_ext           = int(0x8091)
	gl_texture_coord_array_pointer       = int(0x8092)
	gl_texture_coord_array_pointer_ext   = int(0x8092)
	gl_edge_flag_array_pointer           = int(0x8093)
	gl_edge_flag_array_pointer_ext       = int(0x8093)
	gl_interlace_sgix                    = int(0x8094)
	gl_detail_texture_2d_sgis            = int(0x8095)
	gl_detail_texture_2d_binding_sgis    = int(0x8096)
	gl_linear_detail_sgis                = int(0x8097)
	gl_linear_detail_alpha_sgis          = int(0x8098)
	gl_linear_detail_color_sgis          = int(0x8099)
	gl_detail_texture_level_sgis         = int(0x809A)
	gl_detail_texture_mode_sgis          = int(0x809B)
	gl_detail_texture_func_points_sgis   = int(0x809C)
	gl_multisample                       = int(0x809D)
	gl_multisample_arb                   = int(0x809D)
	gl_multisample_ext                   = int(0x809D)
	gl_multisample_sgis                  = int(0x809D)
	gl_sample_alpha_to_coverage          = int(0x809E)
	gl_sample_alpha_to_coverage_arb      = int(0x809E)
	gl_sample_alpha_to_mask_ext          = int(0x809E)
	gl_sample_alpha_to_mask_sgis         = int(0x809E)
	gl_sample_alpha_to_one               = int(0x809F)
	gl_sample_alpha_to_one_arb           = int(0x809F)
	gl_sample_alpha_to_one_ext           = int(0x809F)
	gl_sample_alpha_to_one_sgis          = int(0x809F)
	gl_sample_coverage                   = int(0x80A0)
	gl_sample_coverage_arb               = int(0x80A0)
	gl_sample_mask_ext                   = int(0x80A0)
	gl_sample_mask_sgis                  = int(0x80A0)
	gl_1pass_ext                         = int(0x80A1)
	gl_1pass_sgis                        = int(0x80A1)
	gl_2pass_0_ext                       = int(0x80A2)
	gl_2pass_0_sgis                      = int(0x80A2)
	gl_2pass_1_ext                       = int(0x80A3)
	gl_2pass_1_sgis                      = int(0x80A3)
	gl_4pass_0_ext                       = int(0x80A4)
	gl_4pass_0_sgis                      = int(0x80A4)
	gl_4pass_1_ext                       = int(0x80A5)
	gl_4pass_1_sgis                      = int(0x80A5)
	gl_4pass_2_ext                       = int(0x80A6)
	gl_4pass_2_sgis                      = int(0x80A6)
	gl_4pass_3_ext                       = int(0x80A7)
	gl_4pass_3_sgis                      = int(0x80A7)
	gl_sample_buffers                    = int(0x80A8)
	gl_sample_buffers_arb                = int(0x80A8)
	gl_sample_buffers_ext                = int(0x80A8)
	gl_sample_buffers_sgis               = int(0x80A8)
	gl_samples                           = int(0x80A9)
	gl_samples_arb                       = int(0x80A9)
	gl_samples_ext                       = int(0x80A9)
	gl_samples_sgis                      = int(0x80A9)
	gl_sample_coverage_value             = int(0x80AA)
	gl_sample_coverage_value_arb         = int(0x80AA)
	gl_sample_mask_value_ext             = int(0x80AA)
	gl_sample_mask_value_sgis            = int(0x80AA)
	gl_sample_coverage_invert            = int(0x80AB)
	gl_sample_coverage_invert_arb        = int(0x80AB)
	gl_sample_mask_invert_ext            = int(0x80AB)
	gl_sample_mask_invert_sgis           = int(0x80AB)
	gl_sample_pattern_ext                = int(0x80AC)
	gl_sample_pattern_sgis               = int(0x80AC)
	gl_linear_sharpen_sgis               = int(0x80AD)
	gl_linear_sharpen_alpha_sgis         = int(0x80AE)
	gl_linear_sharpen_color_sgis         = int(0x80AF)
	gl_sharpen_texture_func_points_sgis  = int(0x80B0)
	gl_color_matrix                      = int(0x80B1)
	gl_color_matrix_sgi                  = int(0x80B1)
	gl_color_matrix_stack_depth          = int(0x80B2)
	gl_color_matrix_stack_depth_sgi      = int(0x80B2)
	gl_max_color_matrix_stack_depth      = int(0x80B3)
	gl_max_color_matrix_stack_depth_sgi  = int(0x80B3)
	gl_post_color_matrix_red_scale       = int(0x80B4)
	gl_post_color_matrix_red_scale_sgi   = int(0x80B4)
	gl_post_color_matrix_green_scale     = int(0x80B5)
	gl_post_color_matrix_green_scale_sgi = int(0x80B5)
	gl_post_color_matrix_blue_scale      = int(0x80B6)
	gl_post_color_matrix_blue_scale_sgi  = int(0x80B6)
	gl_post_color_matrix_alpha_scale     = int(0x80B7)
	gl_post_color_matrix_alpha_scale_sgi = int(0x80B7)
	gl_post_color_matrix_red_bias        = int(0x80B8)
	gl_post_color_matrix_red_bias_sgi    = int(0x80B8)
	gl_post_color_matrix_green_bias      = int(0x80B9)
	gl_post_color_matrix_green_bias_sgi  = int(0x80B9)
	gl_post_color_matrix_blue_bias       = int(0x80BA)
	gl_post_color_matrix_blue_bias_sgi   = int(0x80BA)
	gl_post_color_matrix_alpha_bias      = int(0x80BB)
	gl_post_color_matrix_alpha_bias_sgi  = int(0x80BB)
	gl_texture_color_table_sgi           = int(0x80BC)
	gl_proxy_texture_color_table_sgi     = int(0x80BD)
	gl_texture_env_bias_sgix             = int(0x80BE)
	gl_shadow_ambient_sgix               = int(0x80BF)
	gl_texture_compare_fail_value_arb    = int(0x80BF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x80C0" end="0x80CF" vendor="ZiiLabs" |>
pub const (
	gl_blend_dst_rgb       = int(0x80C8)
	gl_blend_dst_rgb_ext   = int(0x80C8)
	gl_blend_dst_rgb_oes   = int(0x80C8)
	gl_blend_src_rgb       = int(0x80C9)
	gl_blend_src_rgb_ext   = int(0x80C9)
	gl_blend_src_rgb_oes   = int(0x80C9)
	gl_blend_dst_alpha     = int(0x80CA)
	gl_blend_dst_alpha_ext = int(0x80CA)
	gl_blend_dst_alpha_oes = int(0x80CA)
	gl_blend_src_alpha     = int(0x80CB)
	gl_blend_src_alpha_ext = int(0x80CB)
	gl_blend_src_alpha_oes = int(0x80CB)
	gl_422_ext             = int(0x80CC)
	gl_422_rev_ext         = int(0x80CD)
	gl_422_average_ext     = int(0x80CE)
	gl_422_rev_average_ext = int(0x80CF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x80D0" end="0x80DF" vendor="SGI" |>
pub const (
	gl_color_table                             = int(0x80D0)
	gl_color_table_sgi                         = int(0x80D0)
	gl_post_convolution_color_table            = int(0x80D1)
	gl_post_convolution_color_table_sgi        = int(0x80D1)
	gl_post_color_matrix_color_table           = int(0x80D2)
	gl_post_color_matrix_color_table_sgi       = int(0x80D2)
	gl_proxy_color_table                       = int(0x80D3)
	gl_proxy_color_table_sgi                   = int(0x80D3)
	gl_proxy_post_convolution_color_table      = int(0x80D4)
	gl_proxy_post_convolution_color_table_sgi  = int(0x80D4)
	gl_proxy_post_color_matrix_color_table     = int(0x80D5)
	gl_proxy_post_color_matrix_color_table_sgi = int(0x80D5)
	gl_color_table_scale                       = int(0x80D6)
	gl_color_table_scale_sgi                   = int(0x80D6)
	gl_color_table_bias                        = int(0x80D7)
	gl_color_table_bias_sgi                    = int(0x80D7)
	gl_color_table_format                      = int(0x80D8)
	gl_color_table_format_sgi                  = int(0x80D8)
	gl_color_table_width                       = int(0x80D9)
	gl_color_table_width_sgi                   = int(0x80D9)
	gl_color_table_red_size                    = int(0x80DA)
	gl_color_table_red_size_sgi                = int(0x80DA)
	gl_color_table_green_size                  = int(0x80DB)
	gl_color_table_green_size_sgi              = int(0x80DB)
	gl_color_table_blue_size                   = int(0x80DC)
	gl_color_table_blue_size_sgi               = int(0x80DC)
	gl_color_table_alpha_size                  = int(0x80DD)
	gl_color_table_alpha_size_sgi              = int(0x80DD)
	gl_color_table_luminance_size              = int(0x80DE)
	gl_color_table_luminance_size_sgi          = int(0x80DE)
	gl_color_table_intensity_size              = int(0x80DF)
	gl_color_table_intensity_size_sgi          = int(0x80DF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x80E0" end="0x810F" vendor="MS" |>
pub const (
	gl_bgr                           = int(0x80E0)
	gl_bgr_ext                       = int(0x80E0)
	gl_bgra                          = int(0x80E1)
	gl_bgra_ext                      = int(0x80E1)
	gl_bgra_img                      = int(0x80E1)
	gl_color_index1_ext              = int(0x80E2)
	gl_color_index2_ext              = int(0x80E3)
	gl_color_index4_ext              = int(0x80E4)
	gl_color_index8_ext              = int(0x80E5)
	gl_color_index12_ext             = int(0x80E6)
	gl_color_index16_ext             = int(0x80E7)
	gl_max_elements_vertices         = int(0x80E8)
	gl_max_elements_vertices_ext     = int(0x80E8)
	gl_max_elements_indices          = int(0x80E9)
	gl_max_elements_indices_ext      = int(0x80E9)
	gl_phong_win                     = int(0x80EA)
	gl_phong_hint_win                = int(0x80EB)
	gl_fog_specular_texture_win      = int(0x80EC)
	gl_texture_index_size_ext        = int(0x80ED)
	gl_parameter_buffer              = int(0x80EE)
	gl_parameter_buffer_arb          = int(0x80EE)
	gl_parameter_buffer_binding      = int(0x80EF)
	gl_parameter_buffer_binding_arb  = int(0x80EF)
	gl_clip_volume_clipping_hint_ext = int(0x80F0)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8110" end="0x814F" vendor="SGI" |>
pub const (
	gl_dual_alpha4_sgis                = int(0x8110)
	gl_dual_alpha8_sgis                = int(0x8111)
	gl_dual_alpha12_sgis               = int(0x8112)
	gl_dual_alpha16_sgis               = int(0x8113)
	gl_dual_luminance4_sgis            = int(0x8114)
	gl_dual_luminance8_sgis            = int(0x8115)
	gl_dual_luminance12_sgis           = int(0x8116)
	gl_dual_luminance16_sgis           = int(0x8117)
	gl_dual_intensity4_sgis            = int(0x8118)
	gl_dual_intensity8_sgis            = int(0x8119)
	gl_dual_intensity12_sgis           = int(0x811A)
	gl_dual_intensity16_sgis           = int(0x811B)
	gl_dual_luminance_alpha4_sgis      = int(0x811C)
	gl_dual_luminance_alpha8_sgis      = int(0x811D)
	gl_quad_alpha4_sgis                = int(0x811E)
	gl_quad_alpha8_sgis                = int(0x811F)
	gl_quad_luminance4_sgis            = int(0x8120)
	gl_quad_luminance8_sgis            = int(0x8121)
	gl_quad_intensity4_sgis            = int(0x8122)
	gl_quad_intensity8_sgis            = int(0x8123)
	gl_dual_texture_select_sgis        = int(0x8124)
	gl_quad_texture_select_sgis        = int(0x8125)
	gl_point_size_min                  = int(0x8126)
	gl_point_size_min_arb              = int(0x8126)
	gl_point_size_min_ext              = int(0x8126)
	gl_point_size_min_sgis             = int(0x8126)
	gl_point_size_max                  = int(0x8127)
	gl_point_size_max_arb              = int(0x8127)
	gl_point_size_max_ext              = int(0x8127)
	gl_point_size_max_sgis             = int(0x8127)
	gl_point_fade_threshold_size       = int(0x8128)
	gl_point_fade_threshold_size_arb   = int(0x8128)
	gl_point_fade_threshold_size_ext   = int(0x8128)
	gl_point_fade_threshold_size_sgis  = int(0x8128)
	gl_distance_attenuation_ext        = int(0x8129)
	gl_distance_attenuation_sgis       = int(0x8129)
	gl_point_distance_attenuation      = int(0x8129)
	gl_point_distance_attenuation_arb  = int(0x8129)
	gl_fog_func_sgis                   = int(0x812A)
	gl_fog_func_points_sgis            = int(0x812B)
	gl_max_fog_func_points_sgis        = int(0x812C)
	gl_clamp_to_border                 = int(0x812D)
	gl_clamp_to_border_arb             = int(0x812D)
	gl_clamp_to_border_ext             = int(0x812D)
	gl_clamp_to_border_nv              = int(0x812D)
	gl_clamp_to_border_sgis            = int(0x812D)
	gl_clamp_to_border_oes             = int(0x812D)
	gl_texture_multi_buffer_hint_sgix  = int(0x812E)
	gl_clamp_to_edge                   = int(0x812F)
	gl_clamp_to_edge_sgis              = int(0x812F)
	gl_pack_skip_volumes_sgis          = int(0x8130)
	gl_pack_image_depth_sgis           = int(0x8131)
	gl_unpack_skip_volumes_sgis        = int(0x8132)
	gl_unpack_image_depth_sgis         = int(0x8133)
	gl_texture_4d_sgis                 = int(0x8134)
	gl_proxy_texture_4d_sgis           = int(0x8135)
	gl_texture_4dsize_sgis             = int(0x8136)
	gl_texture_wrap_q_sgis             = int(0x8137)
	gl_max_4d_texture_size_sgis        = int(0x8138)
	gl_pixel_tex_gen_sgix              = int(0x8139)
	gl_texture_min_lod                 = int(0x813A)
	gl_texture_min_lod_sgis            = int(0x813A)
	gl_texture_max_lod                 = int(0x813B)
	gl_texture_max_lod_sgis            = int(0x813B)
	gl_texture_base_level              = int(0x813C)
	gl_texture_base_level_sgis         = int(0x813C)
	gl_texture_max_level               = int(0x813D)
	gl_texture_max_level_apple         = int(0x813D)
	gl_texture_max_level_sgis          = int(0x813D)
	gl_pixel_tile_best_alignment_sgix  = int(0x813E)
	gl_pixel_tile_cache_increment_sgix = int(0x813F)
	gl_pixel_tile_width_sgix           = int(0x8140)
	gl_pixel_tile_height_sgix          = int(0x8141)
	gl_pixel_tile_grid_width_sgix      = int(0x8142)
	gl_pixel_tile_grid_height_sgix     = int(0x8143)
	gl_pixel_tile_grid_depth_sgix      = int(0x8144)
	gl_pixel_tile_cache_size_sgix      = int(0x8145)
	gl_filter4_sgis                    = int(0x8146)
	gl_texture_filter4_size_sgis       = int(0x8147)
	gl_sprite_sgix                     = int(0x8148)
	gl_sprite_mode_sgix                = int(0x8149)
	gl_sprite_axis_sgix                = int(0x814A)
	gl_sprite_translation_sgix         = int(0x814B)
	gl_sprite_axial_sgix               = int(0x814C)
	gl_sprite_object_aligned_sgix      = int(0x814D)
	gl_sprite_eye_aligned_sgix         = int(0x814E)
	gl_texture_4d_binding_sgis         = int(0x814F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8150" end="0x816F" vendor="HP" |>
pub const (
	gl_ignore_border_hp                          = int(0x8150)
	gl_constant_border                           = int(0x8151)
	gl_constant_border_hp                        = int(0x8151)
	gl_replicate_border                          = int(0x8153)
	gl_replicate_border_hp                       = int(0x8153)
	gl_convolution_border_color                  = int(0x8154)
	gl_convolution_border_color_hp               = int(0x8154)
	gl_image_scale_x_hp                          = int(0x8155)
	gl_image_scale_y_hp                          = int(0x8156)
	gl_image_translate_x_hp                      = int(0x8157)
	gl_image_translate_y_hp                      = int(0x8158)
	gl_image_rotate_angle_hp                     = int(0x8159)
	gl_image_rotate_origin_x_hp                  = int(0x815A)
	gl_image_rotate_origin_y_hp                  = int(0x815B)
	gl_image_mag_filter_hp                       = int(0x815C)
	gl_image_min_filter_hp                       = int(0x815D)
	gl_image_cubic_weight_hp                     = int(0x815E)
	gl_cubic_hp                                  = int(0x815F)
	gl_average_hp                                = int(0x8160)
	gl_image_transform_2d_hp                     = int(0x8161)
	gl_post_image_transform_color_table_hp       = int(0x8162)
	gl_proxy_post_image_transform_color_table_hp = int(0x8163)
	gl_occlusion_test_hp                         = int(0x8165)
	gl_occlusion_test_result_hp                  = int(0x8166)
	gl_texture_lighting_mode_hp                  = int(0x8167)
	gl_texture_post_specular_hp                  = int(0x8168)
	gl_texture_pre_specular_hp                   = int(0x8169)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8170" end="0x81CF" vendor="SGI" |>
pub const (
	gl_linear_clipmap_linear_sgix           = int(0x8170)
	gl_texture_clipmap_center_sgix          = int(0x8171)
	gl_texture_clipmap_frame_sgix           = int(0x8172)
	gl_texture_clipmap_offset_sgix          = int(0x8173)
	gl_texture_clipmap_virtual_depth_sgix   = int(0x8174)
	gl_texture_clipmap_lod_offset_sgix      = int(0x8175)
	gl_texture_clipmap_depth_sgix           = int(0x8176)
	gl_max_clipmap_depth_sgix               = int(0x8177)
	gl_max_clipmap_virtual_depth_sgix       = int(0x8178)
	gl_post_texture_filter_bias_sgix        = int(0x8179)
	gl_post_texture_filter_scale_sgix       = int(0x817A)
	gl_post_texture_filter_bias_range_sgix  = int(0x817B)
	gl_post_texture_filter_scale_range_sgix = int(0x817C)
	gl_reference_plane_sgix                 = int(0x817D)
	gl_reference_plane_equation_sgix        = int(0x817E)
	gl_ir_instrument1_sgix                  = int(0x817F)
	gl_instrument_buffer_pointer_sgix       = int(0x8180)
	gl_instrument_measurements_sgix         = int(0x8181)
	gl_list_priority_sgix                   = int(0x8182)
	gl_calligraphic_fragment_sgix           = int(0x8183)
	gl_pixel_tex_gen_q_ceiling_sgix         = int(0x8184)
	gl_pixel_tex_gen_q_round_sgix           = int(0x8185)
	gl_pixel_tex_gen_q_floor_sgix           = int(0x8186)
	gl_pixel_tex_gen_alpha_ls_sgix          = int(0x8189)
	gl_pixel_tex_gen_alpha_ms_sgix          = int(0x818A)
	gl_framezoom_sgix                       = int(0x818B)
	gl_framezoom_factor_sgix                = int(0x818C)
	gl_max_framezoom_factor_sgix            = int(0x818D)
	gl_texture_lod_bias_s_sgix              = int(0x818E)
	gl_texture_lod_bias_t_sgix              = int(0x818F)
	gl_texture_lod_bias_r_sgix              = int(0x8190)
	gl_generate_mipmap                      = int(0x8191)
	gl_generate_mipmap_sgis                 = int(0x8191)
	gl_generate_mipmap_hint                 = int(0x8192)
	gl_generate_mipmap_hint_sgis            = int(0x8192)
	gl_geometry_deformation_sgix            = int(0x8194)
	gl_texture_deformation_sgix             = int(0x8195)
	gl_deformations_mask_sgix               = int(0x8196)
	gl_max_deformation_order_sgix           = int(0x8197)
	gl_fog_offset_sgix                      = int(0x8198)
	gl_fog_offset_value_sgix                = int(0x8199)
	gl_texture_compare_sgix                 = int(0x819A)
	gl_texture_compare_operator_sgix        = int(0x819B)
	gl_texture_lequal_r_sgix                = int(0x819C)
	gl_texture_gequal_r_sgix                = int(0x819D)
	gl_depth_component16                    = int(0x81A5)
	gl_depth_component16_arb                = int(0x81A5)
	gl_depth_component16_oes                = int(0x81A5)
	gl_depth_component16_sgix               = int(0x81A5)
	gl_depth_component24                    = int(0x81A6)
	gl_depth_component24_arb                = int(0x81A6)
	gl_depth_component24_oes                = int(0x81A6)
	gl_depth_component24_sgix               = int(0x81A6)
	gl_depth_component32                    = int(0x81A7)
	gl_depth_component32_arb                = int(0x81A7)
	gl_depth_component32_oes                = int(0x81A7)
	gl_depth_component32_sgix               = int(0x81A7)
	gl_array_element_lock_first_ext         = int(0x81A8)
	gl_array_element_lock_count_ext         = int(0x81A9)
	gl_cull_vertex_ext                      = int(0x81AA)
	gl_cull_vertex_eye_position_ext         = int(0x81AB)
	gl_cull_vertex_object_position_ext      = int(0x81AC)
	gl_iui_v2f_ext                          = int(0x81AD)
	gl_iui_v3f_ext                          = int(0x81AE)
	gl_iui_n3f_v2f_ext                      = int(0x81AF)
	gl_iui_n3f_v3f_ext                      = int(0x81B0)
	gl_t2f_iui_v2f_ext                      = int(0x81B1)
	gl_t2f_iui_v3f_ext                      = int(0x81B2)
	gl_t2f_iui_n3f_v2f_ext                  = int(0x81B3)
	gl_t2f_iui_n3f_v3f_ext                  = int(0x81B4)
	gl_index_test_ext                       = int(0x81B5)
	gl_index_test_func_ext                  = int(0x81B6)
	gl_index_test_ref_ext                   = int(0x81B7)
	gl_index_material_ext                   = int(0x81B8)
	gl_index_material_parameter_ext         = int(0x81B9)
	gl_index_material_face_ext              = int(0x81BA)
	gl_ycrcb_422_sgix                       = int(0x81BB)
	gl_ycrcb_444_sgix                       = int(0x81BC)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x81D0" end="0x81DF" vendor="SUN" |>
pub const (
	gl_wrap_border_sun            = int(0x81D4)
	gl_unpack_constant_data_sunx  = int(0x81D5)
	gl_texture_constant_data_sunx = int(0x81D6)
	gl_triangle_list_sun          = int(0x81D7)
	gl_replacement_code_sun       = int(0x81D8)
	gl_global_alpha_sun           = int(0x81D9)
	gl_global_alpha_factor_sun    = int(0x81DA)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x81E0" end="0x81FF" vendor="SGI" |>
pub const (
	gl_texture_color_writemask_sgis  = int(0x81EF)
	gl_eye_distance_to_point_sgis    = int(0x81F0)
	gl_object_distance_to_point_sgis = int(0x81F1)
	gl_eye_distance_to_line_sgis     = int(0x81F2)
	gl_object_distance_to_line_sgis  = int(0x81F3)
	gl_eye_point_sgis                = int(0x81F4)
	gl_object_point_sgis             = int(0x81F5)
	gl_eye_line_sgis                 = int(0x81F6)
	gl_object_line_sgis              = int(0x81F7)
	gl_light_model_color_control     = int(0x81F8)
	gl_light_model_color_control_ext = int(0x81F8)
	gl_single_color                  = int(0x81F9)
	gl_single_color_ext              = int(0x81F9)
	gl_separate_specular_color       = int(0x81FA)
	gl_separate_specular_color_ext   = int(0x81FA)
	gl_shared_texture_palette_ext    = int(0x81FB)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8200" end="0x820F" vendor="AMD" comment="Range released by MS 2002/9/16" |>
pub const (
	gl_text_fragment_shader_ati = int(0x8200)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8210" end="0x823F" vendor="ARB" |>
pub const (
	gl_framebuffer_attachment_color_encoding       = int(0x8210)
	gl_framebuffer_attachment_color_encoding_ext   = int(0x8210)
	gl_framebuffer_attachment_component_type       = int(0x8211)
	gl_framebuffer_attachment_component_type_ext   = int(0x8211)
	gl_framebuffer_attachment_red_size             = int(0x8212)
	gl_framebuffer_attachment_green_size           = int(0x8213)
	gl_framebuffer_attachment_blue_size            = int(0x8214)
	gl_framebuffer_attachment_alpha_size           = int(0x8215)
	gl_framebuffer_attachment_depth_size           = int(0x8216)
	gl_framebuffer_attachment_stencil_size         = int(0x8217)
	gl_framebuffer_default                         = int(0x8218)
	gl_framebuffer_undefined                       = int(0x8219)
	gl_framebuffer_undefined_oes                   = int(0x8219)
	gl_depth_stencil_attachment                    = int(0x821A)
	gl_major_version                               = int(0x821B)
	gl_minor_version                               = int(0x821C)
	gl_num_extensions                              = int(0x821D)
	gl_context_flags                               = int(0x821E)
	gl_buffer_immutable_storage                    = int(0x821F)
	gl_buffer_immutable_storage_ext                = int(0x821F)
	gl_buffer_storage_flags                        = int(0x8220)
	gl_buffer_storage_flags_ext                    = int(0x8220)
	gl_primitive_restart_for_patches_supported     = int(0x8221)
	gl_primitive_restart_for_patches_supported_oes = int(0x8221)
	gl_index                                       = int(0x8222)
	gl_compressed_red                              = int(0x8225)
	gl_compressed_rg                               = int(0x8226)
	gl_rg                                          = int(0x8227)
	gl_rg_ext                                      = int(0x8227)
	gl_rg_integer                                  = int(0x8228)
	gl_r8                                          = int(0x8229)
	gl_r8_ext                                      = int(0x8229)
	gl_r16                                         = int(0x822A)
	gl_r16_ext                                     = int(0x822A)
	gl_rg8                                         = int(0x822B)
	gl_rg8_ext                                     = int(0x822B)
	gl_rg16                                        = int(0x822C)
	gl_rg16_ext                                    = int(0x822C)
	gl_r16f                                        = int(0x822D)
	gl_r16f_ext                                    = int(0x822D)
	gl_r32f                                        = int(0x822E)
	gl_r32f_ext                                    = int(0x822E)
	gl_rg16f                                       = int(0x822F)
	gl_rg16f_ext                                   = int(0x822F)
	gl_rg32f                                       = int(0x8230)
	gl_rg32f_ext                                   = int(0x8230)
	gl_r8i                                         = int(0x8231)
	gl_r8ui                                        = int(0x8232)
	gl_r16i                                        = int(0x8233)
	gl_r16ui                                       = int(0x8234)
	gl_r32i                                        = int(0x8235)
	gl_r32ui                                       = int(0x8236)
	gl_rg8i                                        = int(0x8237)
	gl_rg8ui                                       = int(0x8238)
	gl_rg16i                                       = int(0x8239)
	gl_rg16ui                                      = int(0x823A)
	gl_rg32i                                       = int(0x823B)
	gl_rg32ui                                      = int(0x823C)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8240" end="0x82AF" vendor="ARB" comment="Range released by MS on 2002/9/16" |>
pub const (
	gl_sync_cl_event_arb                       = int(0x8240)
	gl_sync_cl_event_complete_arb              = int(0x8241)
	gl_debug_output_synchronous                = int(0x8242)
	gl_debug_output_synchronous_arb            = int(0x8242)
	gl_debug_output_synchronous_khr            = int(0x8242)
	gl_debug_next_logged_message_length        = int(0x8243)
	gl_debug_next_logged_message_length_arb    = int(0x8243)
	gl_debug_next_logged_message_length_khr    = int(0x8243)
	gl_debug_callback_function                 = int(0x8244)
	gl_debug_callback_function_arb             = int(0x8244)
	gl_debug_callback_function_khr             = int(0x8244)
	gl_debug_callback_user_param               = int(0x8245)
	gl_debug_callback_user_param_arb           = int(0x8245)
	gl_debug_callback_user_param_khr           = int(0x8245)
	gl_debug_source_api                        = int(0x8246)
	gl_debug_source_api_arb                    = int(0x8246)
	gl_debug_source_api_khr                    = int(0x8246)
	gl_debug_source_window_system              = int(0x8247)
	gl_debug_source_window_system_arb          = int(0x8247)
	gl_debug_source_window_system_khr          = int(0x8247)
	gl_debug_source_shader_compiler            = int(0x8248)
	gl_debug_source_shader_compiler_arb        = int(0x8248)
	gl_debug_source_shader_compiler_khr        = int(0x8248)
	gl_debug_source_third_party                = int(0x8249)
	gl_debug_source_third_party_arb            = int(0x8249)
	gl_debug_source_third_party_khr            = int(0x8249)
	gl_debug_source_application                = int(0x824A)
	gl_debug_source_application_arb            = int(0x824A)
	gl_debug_source_application_khr            = int(0x824A)
	gl_debug_source_other                      = int(0x824B)
	gl_debug_source_other_arb                  = int(0x824B)
	gl_debug_source_other_khr                  = int(0x824B)
	gl_debug_type_error                        = int(0x824C)
	gl_debug_type_error_arb                    = int(0x824C)
	gl_debug_type_error_khr                    = int(0x824C)
	gl_debug_type_deprecated_behavior          = int(0x824D)
	gl_debug_type_deprecated_behavior_arb      = int(0x824D)
	gl_debug_type_deprecated_behavior_khr      = int(0x824D)
	gl_debug_type_undefined_behavior           = int(0x824E)
	gl_debug_type_undefined_behavior_arb       = int(0x824E)
	gl_debug_type_undefined_behavior_khr       = int(0x824E)
	gl_debug_type_portability                  = int(0x824F)
	gl_debug_type_portability_arb              = int(0x824F)
	gl_debug_type_portability_khr              = int(0x824F)
	gl_debug_type_performance                  = int(0x8250)
	gl_debug_type_performance_arb              = int(0x8250)
	gl_debug_type_performance_khr              = int(0x8250)
	gl_debug_type_other                        = int(0x8251)
	gl_debug_type_other_arb                    = int(0x8251)
	gl_debug_type_other_khr                    = int(0x8251)
	gl_lose_context_on_reset                   = int(0x8252)
	gl_lose_context_on_reset_arb               = int(0x8252)
	gl_lose_context_on_reset_ext               = int(0x8252)
	gl_lose_context_on_reset_khr               = int(0x8252)
	gl_guilty_context_reset                    = int(0x8253)
	gl_guilty_context_reset_arb                = int(0x8253)
	gl_guilty_context_reset_ext                = int(0x8253)
	gl_guilty_context_reset_khr                = int(0x8253)
	gl_innocent_context_reset                  = int(0x8254)
	gl_innocent_context_reset_arb              = int(0x8254)
	gl_innocent_context_reset_ext              = int(0x8254)
	gl_innocent_context_reset_khr              = int(0x8254)
	gl_unknown_context_reset                   = int(0x8255)
	gl_unknown_context_reset_arb               = int(0x8255)
	gl_unknown_context_reset_ext               = int(0x8255)
	gl_unknown_context_reset_khr               = int(0x8255)
	gl_reset_notification_strategy             = int(0x8256)
	gl_reset_notification_strategy_arb         = int(0x8256)
	gl_reset_notification_strategy_ext         = int(0x8256)
	gl_reset_notification_strategy_khr         = int(0x8256)
	gl_program_binary_retrievable_hint         = int(0x8257)
	gl_program_separable                       = int(0x8258)
	gl_program_separable_ext                   = int(0x8258)
	gl_active_program                          = int(0x8259)
	gl_active_program_ext                      = int(0x8259)
	gl_program_pipeline_binding                = int(0x825A)
	gl_program_pipeline_binding_ext            = int(0x825A)
	gl_max_viewports                           = int(0x825B)
	gl_max_viewports_nv                        = int(0x825B)
	gl_max_viewports_oes                       = int(0x825B)
	gl_viewport_subpixel_bits                  = int(0x825C)
	gl_viewport_subpixel_bits_ext              = int(0x825C)
	gl_viewport_subpixel_bits_nv               = int(0x825C)
	gl_viewport_subpixel_bits_oes              = int(0x825C)
	gl_viewport_bounds_range                   = int(0x825D)
	gl_viewport_bounds_range_ext               = int(0x825D)
	gl_viewport_bounds_range_nv                = int(0x825D)
	gl_viewport_bounds_range_oes               = int(0x825D)
	gl_layer_provoking_vertex                  = int(0x825E)
	gl_layer_provoking_vertex_ext              = int(0x825E)
	gl_layer_provoking_vertex_oes              = int(0x825E)
	gl_viewport_index_provoking_vertex         = int(0x825F)
	gl_viewport_index_provoking_vertex_ext     = int(0x825F)
	gl_viewport_index_provoking_vertex_nv      = int(0x825F)
	gl_viewport_index_provoking_vertex_oes     = int(0x825F)
	gl_undefined_vertex                        = int(0x8260)
	gl_undefined_vertex_ext                    = int(0x8260)
	gl_undefined_vertex_oes                    = int(0x8260)
	gl_no_reset_notification                   = int(0x8261)
	gl_no_reset_notification_arb               = int(0x8261)
	gl_no_reset_notification_ext               = int(0x8261)
	gl_no_reset_notification_khr               = int(0x8261)
	gl_max_compute_shared_memory_size          = int(0x8262)
	gl_max_compute_uniform_components          = int(0x8263)
	gl_max_compute_atomic_counter_buffers      = int(0x8264)
	gl_max_compute_atomic_counters             = int(0x8265)
	gl_max_combined_compute_uniform_components = int(0x8266)
	gl_compute_work_group_size                 = int(0x8267)
	gl_debug_type_marker                       = int(0x8268)
	gl_debug_type_marker_khr                   = int(0x8268)
	gl_debug_type_push_group                   = int(0x8269)
	gl_debug_type_push_group_khr               = int(0x8269)
	gl_debug_type_pop_group                    = int(0x826A)
	gl_debug_type_pop_group_khr                = int(0x826A)
	gl_debug_severity_notification             = int(0x826B)
	gl_debug_severity_notification_khr         = int(0x826B)
	gl_max_debug_group_stack_depth             = int(0x826C)
	gl_max_debug_group_stack_depth_khr         = int(0x826C)
	gl_debug_group_stack_depth                 = int(0x826D)
	gl_debug_group_stack_depth_khr             = int(0x826D)
	gl_max_uniform_locations                   = int(0x826E)
	gl_internalformat_supported                = int(0x826F)
	gl_internalformat_preferred                = int(0x8270)
	gl_internalformat_red_size                 = int(0x8271)
	gl_internalformat_green_size               = int(0x8272)
	gl_internalformat_blue_size                = int(0x8273)
	gl_internalformat_alpha_size               = int(0x8274)
	gl_internalformat_depth_size               = int(0x8275)
	gl_internalformat_stencil_size             = int(0x8276)
	gl_internalformat_shared_size              = int(0x8277)
	gl_internalformat_red_type                 = int(0x8278)
	gl_internalformat_green_type               = int(0x8279)
	gl_internalformat_blue_type                = int(0x827A)
	gl_internalformat_alpha_type               = int(0x827B)
	gl_internalformat_depth_type               = int(0x827C)
	gl_internalformat_stencil_type             = int(0x827D)
	gl_max_width                               = int(0x827E)
	gl_max_height                              = int(0x827F)
	gl_max_depth                               = int(0x8280)
	gl_max_layers                              = int(0x8281)
	gl_max_combined_dimensions                 = int(0x8282)
	gl_color_components                        = int(0x8283)
	gl_depth_components                        = int(0x8284)
	gl_stencil_components                      = int(0x8285)
	gl_color_renderable                        = int(0x8286)
	gl_depth_renderable                        = int(0x8287)
	gl_stencil_renderable                      = int(0x8288)
	gl_framebuffer_renderable                  = int(0x8289)
	gl_framebuffer_renderable_layered          = int(0x828A)
	gl_framebuffer_blend                       = int(0x828B)
	gl_read_pixels                             = int(0x828C)
	gl_read_pixels_format                      = int(0x828D)
	gl_read_pixels_type                        = int(0x828E)
	gl_texture_image_format                    = int(0x828F)
	gl_texture_image_type                      = int(0x8290)
	gl_get_texture_image_format                = int(0x8291)
	gl_get_texture_image_type                  = int(0x8292)
	gl_mipmap                                  = int(0x8293)
	gl_manual_generate_mipmap                  = int(0x8294)
	gl_auto_generate_mipmap                    = int(0x8295)
	gl_color_encoding                          = int(0x8296)
	gl_srgb_read                               = int(0x8297)
	gl_srgb_write                              = int(0x8298)
	gl_srgb_decode_arb                         = int(0x8299)
	gl_filter                                  = int(0x829A)
	gl_vertex_texture                          = int(0x829B)
	gl_tess_control_texture                    = int(0x829C)
	gl_tess_evaluation_texture                 = int(0x829D)
	gl_geometry_texture                        = int(0x829E)
	gl_fragment_texture                        = int(0x829F)
	gl_compute_texture                         = int(0x82A0)
	gl_texture_shadow                          = int(0x82A1)
	gl_texture_gather                          = int(0x82A2)
	gl_texture_gather_shadow                   = int(0x82A3)
	gl_shader_image_load                       = int(0x82A4)
	gl_shader_image_store                      = int(0x82A5)
	gl_shader_image_atomic                     = int(0x82A6)
	gl_image_texel_size                        = int(0x82A7)
	gl_image_compatibility_class               = int(0x82A8)
	gl_image_pixel_format                      = int(0x82A9)
	gl_image_pixel_type                        = int(0x82AA)
	gl_simultaneous_texture_and_depth_test     = int(0x82AC)
	gl_simultaneous_texture_and_stencil_test   = int(0x82AD)
	gl_simultaneous_texture_and_depth_write    = int(0x82AE)
	gl_simultaneous_texture_and_stencil_write  = int(0x82AF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x82B0" end="0x830F" vendor="ARB" comment="Range reclaimed from ADD on 2012/05/10" |>
pub const (
	gl_texture_compressed_block_width           = int(0x82B1)
	gl_texture_compressed_block_height          = int(0x82B2)
	gl_texture_compressed_block_size            = int(0x82B3)
	gl_clear_buffer                             = int(0x82B4)
	gl_texture_view                             = int(0x82B5)
	gl_view_compatibility_class                 = int(0x82B6)
	gl_full_support                             = int(0x82B7)
	gl_caveat_support                           = int(0x82B8)
	gl_image_class_4_x_32                       = int(0x82B9)
	gl_image_class_2_x_32                       = int(0x82BA)
	gl_image_class_1_x_32                       = int(0x82BB)
	gl_image_class_4_x_16                       = int(0x82BC)
	gl_image_class_2_x_16                       = int(0x82BD)
	gl_image_class_1_x_16                       = int(0x82BE)
	gl_image_class_4_x_8                        = int(0x82BF)
	gl_image_class_2_x_8                        = int(0x82C0)
	gl_image_class_1_x_8                        = int(0x82C1)
	gl_image_class_11_11_10                     = int(0x82C2)
	gl_image_class_10_10_10_2                   = int(0x82C3)
	gl_view_class_128_bits                      = int(0x82C4)
	gl_view_class_96_bits                       = int(0x82C5)
	gl_view_class_64_bits                       = int(0x82C6)
	gl_view_class_48_bits                       = int(0x82C7)
	gl_view_class_32_bits                       = int(0x82C8)
	gl_view_class_24_bits                       = int(0x82C9)
	gl_view_class_16_bits                       = int(0x82CA)
	gl_view_class_8_bits                        = int(0x82CB)
	gl_view_class_s3tc_dxt1_rgb                 = int(0x82CC)
	gl_view_class_s3tc_dxt1_rgba                = int(0x82CD)
	gl_view_class_s3tc_dxt3_rgba                = int(0x82CE)
	gl_view_class_s3tc_dxt5_rgba                = int(0x82CF)
	gl_view_class_rgtc1_red                     = int(0x82D0)
	gl_view_class_rgtc2_rg                      = int(0x82D1)
	gl_view_class_bptc_unorm                    = int(0x82D2)
	gl_view_class_bptc_float                    = int(0x82D3)
	gl_vertex_attrib_binding                    = int(0x82D4)
	gl_vertex_attrib_relative_offset            = int(0x82D5)
	gl_vertex_binding_divisor                   = int(0x82D6)
	gl_vertex_binding_offset                    = int(0x82D7)
	gl_vertex_binding_stride                    = int(0x82D8)
	gl_max_vertex_attrib_relative_offset        = int(0x82D9)
	gl_max_vertex_attrib_bindings               = int(0x82DA)
	gl_texture_view_min_level                   = int(0x82DB)
	gl_texture_view_min_level_ext               = int(0x82DB)
	gl_texture_view_min_level_oes               = int(0x82DB)
	gl_texture_view_num_levels                  = int(0x82DC)
	gl_texture_view_num_levels_ext              = int(0x82DC)
	gl_texture_view_num_levels_oes              = int(0x82DC)
	gl_texture_view_min_layer                   = int(0x82DD)
	gl_texture_view_min_layer_ext               = int(0x82DD)
	gl_texture_view_min_layer_oes               = int(0x82DD)
	gl_texture_view_num_layers                  = int(0x82DE)
	gl_texture_view_num_layers_ext              = int(0x82DE)
	gl_texture_view_num_layers_oes              = int(0x82DE)
	gl_texture_immutable_levels                 = int(0x82DF)
	gl_buffer                                   = int(0x82E0)
	gl_buffer_khr                               = int(0x82E0)
	gl_shader                                   = int(0x82E1)
	gl_shader_khr                               = int(0x82E1)
	gl_program                                  = int(0x82E2)
	gl_program_khr                              = int(0x82E2)
	gl_query                                    = int(0x82E3)
	gl_query_khr                                = int(0x82E3)
	gl_program_pipeline                         = int(0x82E4)
	gl_program_pipeline_khr                     = int(0x82E4)
	gl_max_vertex_attrib_stride                 = int(0x82E5)
	gl_sampler                                  = int(0x82E6)
	gl_sampler_khr                              = int(0x82E6)
	gl_display_list                             = int(0x82E7)
	gl_max_label_length                         = int(0x82E8)
	gl_max_label_length_khr                     = int(0x82E8)
	gl_num_shading_language_versions            = int(0x82E9)
	gl_query_target                             = int(0x82EA)
	gl_transform_feedback_overflow              = int(0x82EC)
	gl_transform_feedback_overflow_arb          = int(0x82EC)
	gl_transform_feedback_stream_overflow       = int(0x82ED)
	gl_transform_feedback_stream_overflow_arb   = int(0x82ED)
	gl_vertices_submitted                       = int(0x82EE)
	gl_vertices_submitted_arb                   = int(0x82EE)
	gl_primitives_submitted                     = int(0x82EF)
	gl_primitives_submitted_arb                 = int(0x82EF)
	gl_vertex_shader_invocations                = int(0x82F0)
	gl_vertex_shader_invocations_arb            = int(0x82F0)
	gl_tess_control_shader_patches              = int(0x82F1)
	gl_tess_control_shader_patches_arb          = int(0x82F1)
	gl_tess_evaluation_shader_invocations       = int(0x82F2)
	gl_tess_evaluation_shader_invocations_arb   = int(0x82F2)
	gl_geometry_shader_primitives_emitted       = int(0x82F3)
	gl_geometry_shader_primitives_emitted_arb   = int(0x82F3)
	gl_fragment_shader_invocations              = int(0x82F4)
	gl_fragment_shader_invocations_arb          = int(0x82F4)
	gl_compute_shader_invocations               = int(0x82F5)
	gl_compute_shader_invocations_arb           = int(0x82F5)
	gl_clipping_input_primitives                = int(0x82F6)
	gl_clipping_input_primitives_arb            = int(0x82F6)
	gl_clipping_output_primitives               = int(0x82F7)
	gl_clipping_output_primitives_arb           = int(0x82F7)
	gl_sparse_buffer_page_size_arb              = int(0x82F8)
	gl_max_cull_distances                       = int(0x82F9)
	gl_max_cull_distances_ext                   = int(0x82F9)
	gl_max_combined_clip_and_cull_distances     = int(0x82FA)
	gl_max_combined_clip_and_cull_distances_ext = int(0x82FA)
	gl_context_release_behavior                 = int(0x82FB)
	gl_context_release_behavior_khr             = int(0x82FB)
	gl_context_release_behavior_flush           = int(0x82FC)
	gl_context_release_behavior_flush_khr       = int(0x82FC)
	gl_robust_gpu_timeout_ms_khr                = int(0x82FD)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8310" end="0x832F" vendor="SGI" |>
pub const (
	gl_depth_pass_instrument_sgix          = int(0x8310)
	gl_depth_pass_instrument_counters_sgix = int(0x8311)
	gl_depth_pass_instrument_max_sgix      = int(0x8312)
	gl_fragments_instrument_sgix           = int(0x8313)
	gl_fragments_instrument_counters_sgix  = int(0x8314)
	gl_fragments_instrument_max_sgix       = int(0x8315)
	gl_convolution_hint_sgix               = int(0x8316)
	gl_ycrcb_sgix                          = int(0x8318)
	gl_ycrcba_sgix                         = int(0x8319)
	gl_unpack_compressed_size_sgix         = int(0x831A)
	gl_pack_max_compressed_size_sgix       = int(0x831B)
	gl_pack_compressed_size_sgix           = int(0x831C)
	gl_slim8u_sgix                         = int(0x831D)
	gl_slim10u_sgix                        = int(0x831E)
	gl_slim12s_sgix                        = int(0x831F)
	gl_alpha_min_sgix                      = int(0x8320)
	gl_alpha_max_sgix                      = int(0x8321)
	gl_scalebias_hint_sgix                 = int(0x8322)
	gl_async_marker_sgix                   = int(0x8329)
	gl_pixel_tex_gen_mode_sgix             = int(0x832B)
	gl_async_histogram_sgix                = int(0x832C)
	gl_max_async_histogram_sgix            = int(0x832D)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8330" end="0x833F" vendor="SUN" |>
pub const (
	gl_pixel_transform_2d_ext                 = int(0x8330)
	gl_pixel_mag_filter_ext                   = int(0x8331)
	gl_pixel_min_filter_ext                   = int(0x8332)
	gl_pixel_cubic_weight_ext                 = int(0x8333)
	gl_cubic_ext                              = int(0x8334)
	gl_average_ext                            = int(0x8335)
	gl_pixel_transform_2d_stack_depth_ext     = int(0x8336)
	gl_max_pixel_transform_2d_stack_depth_ext = int(0x8337)
	gl_pixel_transform_2d_matrix_ext          = int(0x8338)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8340" end="0x836F" vendor="SGI" |>
pub const (
	gl_fragment_material_ext            = int(0x8349)
	gl_fragment_normal_ext              = int(0x834A)
	gl_fragment_color_ext               = int(0x834C)
	gl_attenuation_ext                  = int(0x834D)
	gl_shadow_attenuation_ext           = int(0x834E)
	gl_texture_application_mode_ext     = int(0x834F)
	gl_texture_light_ext                = int(0x8350)
	gl_texture_material_face_ext        = int(0x8351)
	gl_texture_material_parameter_ext   = int(0x8352)
	gl_pixel_texture_sgis               = int(0x8353)
	gl_pixel_fragment_rgb_source_sgis   = int(0x8354)
	gl_pixel_fragment_alpha_source_sgis = int(0x8355)
	gl_pixel_group_color_sgis           = int(0x8356)
	gl_line_quality_hint_sgix           = int(0x835B)
	gl_async_tex_image_sgix             = int(0x835C)
	gl_async_draw_pixels_sgix           = int(0x835D)
	gl_async_read_pixels_sgix           = int(0x835E)
	gl_max_async_tex_image_sgix         = int(0x835F)
	gl_max_async_draw_pixels_sgix       = int(0x8360)
	gl_max_async_read_pixels_sgix       = int(0x8361)
	gl_unsigned_byte_2_3_3_rev          = int(0x8362)
	gl_unsigned_byte_2_3_3_rev_ext      = int(0x8362)
	gl_unsigned_short_5_6_5             = int(0x8363)
	gl_unsigned_short_5_6_5_ext         = int(0x8363)
	gl_unsigned_short_5_6_5_rev         = int(0x8364)
	gl_unsigned_short_5_6_5_rev_ext     = int(0x8364)
	gl_unsigned_short_4_4_4_4_rev       = int(0x8365)
	gl_unsigned_short_4_4_4_4_rev_ext   = int(0x8365)
	gl_unsigned_short_4_4_4_4_rev_img   = int(0x8365)
	gl_unsigned_short_1_5_5_5_rev       = int(0x8366)
	gl_unsigned_short_1_5_5_5_rev_ext   = int(0x8366)
	gl_unsigned_int_8_8_8_8_rev         = int(0x8367)
	gl_unsigned_int_8_8_8_8_rev_ext     = int(0x8367)
	gl_unsigned_int_2_10_10_10_rev      = int(0x8368)
	gl_unsigned_int_2_10_10_10_rev_ext  = int(0x8368)
	gl_texture_max_clamp_s_sgix         = int(0x8369)
	gl_texture_max_clamp_t_sgix         = int(0x836A)
	gl_texture_max_clamp_r_sgix         = int(0x836B)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8370" end="0x837F" vendor="HP" |>
pub const (
	gl_mirrored_repeat     = int(0x8370)
	gl_mirrored_repeat_arb = int(0x8370)
	gl_mirrored_repeat_ibm = int(0x8370)
	gl_mirrored_repeat_oes = int(0x8370)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x83A0" end="0x83BF" vendor="S3" |>
pub const (
	gl_rgb_s3tc        = int(0x83A0)
	gl_rgb4_s3tc       = int(0x83A1)
	gl_rgba_s3tc       = int(0x83A2)
	gl_rgba4_s3tc      = int(0x83A3)
	gl_rgba_dxt5_s3tc  = int(0x83A4)
	gl_rgba4_dxt5_s3tc = int(0x83A5)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x83C0" end="0x83EF" vendor="SGI" comment="Most of this could be reclaimed" |>
pub const (
	gl_vertex_preclip_sgix      = int(0x83EE)
	gl_vertex_preclip_hint_sgix = int(0x83EF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x83F0" end="0x83FF" vendor="INTEL" |>
pub const (
	gl_compressed_rgb_s3tc_dxt1_ext                = int(0x83F0)
	gl_compressed_rgba_s3tc_dxt1_ext               = int(0x83F1)
	gl_compressed_rgba_s3tc_dxt3_angle             = int(0x83F2)
	gl_compressed_rgba_s3tc_dxt3_ext               = int(0x83F2)
	gl_compressed_rgba_s3tc_dxt5_angle             = int(0x83F3)
	gl_compressed_rgba_s3tc_dxt5_ext               = int(0x83F3)
	gl_parallel_arrays_intel                       = int(0x83F4)
	gl_vertex_array_parallel_pointers_intel        = int(0x83F5)
	gl_normal_array_parallel_pointers_intel        = int(0x83F6)
	gl_color_array_parallel_pointers_intel         = int(0x83F7)
	gl_texture_coord_array_parallel_pointers_intel = int(0x83F8)
	gl_perfquery_donot_flush_intel                 = int(0x83F9)
	gl_perfquery_flush_intel                       = int(0x83FA)
	gl_perfquery_wait_intel                        = int(0x83FB)
	gl_blackhole_render_intel                      = int(0x83FC)
	gl_conservative_rasterization_intel            = int(0x83FE)
	gl_texture_memory_layout_intel                 = int(0x83FF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8400" end="0x846F" vendor="SGI" |>
pub const (
	gl_fragment_lighting_sgix                         = int(0x8400)
	gl_fragment_color_material_sgix                   = int(0x8401)
	gl_fragment_color_material_face_sgix              = int(0x8402)
	gl_fragment_color_material_parameter_sgix         = int(0x8403)
	gl_max_fragment_lights_sgix                       = int(0x8404)
	gl_max_active_lights_sgix                         = int(0x8405)
	gl_current_raster_normal_sgix                     = int(0x8406)
	gl_light_env_mode_sgix                            = int(0x8407)
	gl_fragment_light_model_local_viewer_sgix         = int(0x8408)
	gl_fragment_light_model_two_side_sgix             = int(0x8409)
	gl_fragment_light_model_ambient_sgix              = int(0x840A)
	gl_fragment_light_model_normal_interpolation_sgix = int(0x840B)
	gl_fragment_light0_sgix                           = int(0x840C)
	gl_fragment_light1_sgix                           = int(0x840D)
	gl_fragment_light2_sgix                           = int(0x840E)
	gl_fragment_light3_sgix                           = int(0x840F)
	gl_fragment_light4_sgix                           = int(0x8410)
	gl_fragment_light5_sgix                           = int(0x8411)
	gl_fragment_light6_sgix                           = int(0x8412)
	gl_fragment_light7_sgix                           = int(0x8413)
	gl_pack_resample_sgix                             = int(0x842E)
	gl_unpack_resample_sgix                           = int(0x842F)
	gl_resample_decimate_sgix                         = int(0x8430)
	gl_resample_replicate_sgix                        = int(0x8433)
	gl_resample_zero_fill_sgix                        = int(0x8434)
	gl_tangent_array_ext                              = int(0x8439)
	gl_binormal_array_ext                             = int(0x843A)
	gl_current_tangent_ext                            = int(0x843B)
	gl_current_binormal_ext                           = int(0x843C)
	gl_tangent_array_type_ext                         = int(0x843E)
	gl_tangent_array_stride_ext                       = int(0x843F)
	gl_binormal_array_type_ext                        = int(0x8440)
	gl_binormal_array_stride_ext                      = int(0x8441)
	gl_tangent_array_pointer_ext                      = int(0x8442)
	gl_binormal_array_pointer_ext                     = int(0x8443)
	gl_map1_tangent_ext                               = int(0x8444)
	gl_map2_tangent_ext                               = int(0x8445)
	gl_map1_binormal_ext                              = int(0x8446)
	gl_map2_binormal_ext                              = int(0x8447)
	gl_nearest_clipmap_nearest_sgix                   = int(0x844D)
	gl_nearest_clipmap_linear_sgix                    = int(0x844E)
	gl_linear_clipmap_nearest_sgix                    = int(0x844F)
	gl_fog_coordinate_source                          = int(0x8450)
	gl_fog_coordinate_source_ext                      = int(0x8450)
	gl_fog_coord_src                                  = int(0x8450)
	gl_fog_coordinate                                 = int(0x8451)
	gl_fog_coordinate_ext                             = int(0x8451)
	gl_fog_coord                                      = int(0x8451)
	gl_fragment_depth                                 = int(0x8452)
	gl_fragment_depth_ext                             = int(0x8452)
	gl_current_fog_coordinate                         = int(0x8453)
	gl_current_fog_coord                              = int(0x8453)
	gl_current_fog_coordinate_ext                     = int(0x8453)
	gl_fog_coordinate_array_type                      = int(0x8454)
	gl_fog_coordinate_array_type_ext                  = int(0x8454)
	gl_fog_coord_array_type                           = int(0x8454)
	gl_fog_coordinate_array_stride                    = int(0x8455)
	gl_fog_coordinate_array_stride_ext                = int(0x8455)
	gl_fog_coord_array_stride                         = int(0x8455)
	gl_fog_coordinate_array_pointer                   = int(0x8456)
	gl_fog_coordinate_array_pointer_ext               = int(0x8456)
	gl_fog_coord_array_pointer                        = int(0x8456)
	gl_fog_coordinate_array                           = int(0x8457)
	gl_fog_coordinate_array_ext                       = int(0x8457)
	gl_fog_coord_array                                = int(0x8457)
	gl_color_sum                                      = int(0x8458)
	gl_color_sum_arb                                  = int(0x8458)
	gl_color_sum_ext                                  = int(0x8458)
	gl_current_secondary_color                        = int(0x8459)
	gl_current_secondary_color_ext                    = int(0x8459)
	gl_secondary_color_array_size                     = int(0x845A)
	gl_secondary_color_array_size_ext                 = int(0x845A)
	gl_secondary_color_array_type                     = int(0x845B)
	gl_secondary_color_array_type_ext                 = int(0x845B)
	gl_secondary_color_array_stride                   = int(0x845C)
	gl_secondary_color_array_stride_ext               = int(0x845C)
	gl_secondary_color_array_pointer                  = int(0x845D)
	gl_secondary_color_array_pointer_ext              = int(0x845D)
	gl_secondary_color_array                          = int(0x845E)
	gl_secondary_color_array_ext                      = int(0x845E)
	gl_current_raster_secondary_color                 = int(0x845F)
	gl_aliased_point_size_range                       = int(0x846D)
	gl_aliased_line_width_range                       = int(0x846E)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8490" end="0x849F" vendor="REND" |>
pub const (
	gl_screen_coordinates_rend = int(0x8490)
	gl_inverted_screen_w_rend  = int(0x8491)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x84C0" end="0x84EF" vendor="ARB" |>
pub const (
	gl_texture0                            = int(0x84C0)
	gl_texture0_arb                        = int(0x84C0)
	gl_texture1                            = int(0x84C1)
	gl_texture1_arb                        = int(0x84C1)
	gl_texture2                            = int(0x84C2)
	gl_texture2_arb                        = int(0x84C2)
	gl_texture3                            = int(0x84C3)
	gl_texture3_arb                        = int(0x84C3)
	gl_texture4                            = int(0x84C4)
	gl_texture4_arb                        = int(0x84C4)
	gl_texture5                            = int(0x84C5)
	gl_texture5_arb                        = int(0x84C5)
	gl_texture6                            = int(0x84C6)
	gl_texture6_arb                        = int(0x84C6)
	gl_texture7                            = int(0x84C7)
	gl_texture7_arb                        = int(0x84C7)
	gl_texture8                            = int(0x84C8)
	gl_texture8_arb                        = int(0x84C8)
	gl_texture9                            = int(0x84C9)
	gl_texture9_arb                        = int(0x84C9)
	gl_texture10                           = int(0x84CA)
	gl_texture10_arb                       = int(0x84CA)
	gl_texture11                           = int(0x84CB)
	gl_texture11_arb                       = int(0x84CB)
	gl_texture12                           = int(0x84CC)
	gl_texture12_arb                       = int(0x84CC)
	gl_texture13                           = int(0x84CD)
	gl_texture13_arb                       = int(0x84CD)
	gl_texture14                           = int(0x84CE)
	gl_texture14_arb                       = int(0x84CE)
	gl_texture15                           = int(0x84CF)
	gl_texture15_arb                       = int(0x84CF)
	gl_texture16                           = int(0x84D0)
	gl_texture16_arb                       = int(0x84D0)
	gl_texture17                           = int(0x84D1)
	gl_texture17_arb                       = int(0x84D1)
	gl_texture18                           = int(0x84D2)
	gl_texture18_arb                       = int(0x84D2)
	gl_texture19                           = int(0x84D3)
	gl_texture19_arb                       = int(0x84D3)
	gl_texture20                           = int(0x84D4)
	gl_texture20_arb                       = int(0x84D4)
	gl_texture21                           = int(0x84D5)
	gl_texture21_arb                       = int(0x84D5)
	gl_texture22                           = int(0x84D6)
	gl_texture22_arb                       = int(0x84D6)
	gl_texture23                           = int(0x84D7)
	gl_texture23_arb                       = int(0x84D7)
	gl_texture24                           = int(0x84D8)
	gl_texture24_arb                       = int(0x84D8)
	gl_texture25                           = int(0x84D9)
	gl_texture25_arb                       = int(0x84D9)
	gl_texture26                           = int(0x84DA)
	gl_texture26_arb                       = int(0x84DA)
	gl_texture27                           = int(0x84DB)
	gl_texture27_arb                       = int(0x84DB)
	gl_texture28                           = int(0x84DC)
	gl_texture28_arb                       = int(0x84DC)
	gl_texture29                           = int(0x84DD)
	gl_texture29_arb                       = int(0x84DD)
	gl_texture30                           = int(0x84DE)
	gl_texture30_arb                       = int(0x84DE)
	gl_texture31                           = int(0x84DF)
	gl_texture31_arb                       = int(0x84DF)
	gl_active_texture                      = int(0x84E0)
	gl_active_texture_arb                  = int(0x84E0)
	gl_client_active_texture               = int(0x84E1)
	gl_client_active_texture_arb           = int(0x84E1)
	gl_max_texture_units                   = int(0x84E2)
	gl_max_texture_units_arb               = int(0x84E2)
	gl_transpose_modelview_matrix          = int(0x84E3)
	gl_transpose_modelview_matrix_arb      = int(0x84E3)
	gl_path_transpose_modelview_matrix_nv  = int(0x84E3)
	gl_transpose_projection_matrix         = int(0x84E4)
	gl_transpose_projection_matrix_arb     = int(0x84E4)
	gl_path_transpose_projection_matrix_nv = int(0x84E4)
	gl_transpose_texture_matrix            = int(0x84E5)
	gl_transpose_texture_matrix_arb        = int(0x84E5)
	gl_transpose_color_matrix              = int(0x84E6)
	gl_transpose_color_matrix_arb          = int(0x84E6)
	gl_subtract                            = int(0x84E7)
	gl_subtract_arb                        = int(0x84E7)
	gl_max_renderbuffer_size               = int(0x84E8)
	gl_max_renderbuffer_size_ext           = int(0x84E8)
	gl_max_renderbuffer_size_oes           = int(0x84E8)
	gl_compressed_alpha                    = int(0x84E9)
	gl_compressed_alpha_arb                = int(0x84E9)
	gl_compressed_luminance                = int(0x84EA)
	gl_compressed_luminance_arb            = int(0x84EA)
	gl_compressed_luminance_alpha          = int(0x84EB)
	gl_compressed_luminance_alpha_arb      = int(0x84EB)
	gl_compressed_intensity                = int(0x84EC)
	gl_compressed_intensity_arb            = int(0x84EC)
	gl_compressed_rgb                      = int(0x84ED)
	gl_compressed_rgb_arb                  = int(0x84ED)
	gl_compressed_rgba                     = int(0x84EE)
	gl_compressed_rgba_arb                 = int(0x84EE)
	gl_texture_compression_hint            = int(0x84EF)
	gl_texture_compression_hint_arb        = int(0x84EF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x84F0" end="0x855F" vendor="NV" |>
pub const (
	gl_uniform_block_referenced_by_tess_control_shader    = int(0x84F0)
	gl_uniform_block_referenced_by_tess_evaluation_shader = int(0x84F1)
	gl_all_completed_nv                                   = int(0x84F2)
	gl_fence_status_nv                                    = int(0x84F3)
	gl_fence_condition_nv                                 = int(0x84F4)
	gl_texture_rectangle                                  = int(0x84F5)
	gl_texture_rectangle_arb                              = int(0x84F5)
	gl_texture_rectangle_nv                               = int(0x84F5)
	gl_texture_binding_rectangle                          = int(0x84F6)
	gl_texture_binding_rectangle_arb                      = int(0x84F6)
	gl_texture_binding_rectangle_nv                       = int(0x84F6)
	gl_proxy_texture_rectangle                            = int(0x84F7)
	gl_proxy_texture_rectangle_arb                        = int(0x84F7)
	gl_proxy_texture_rectangle_nv                         = int(0x84F7)
	gl_max_rectangle_texture_size                         = int(0x84F8)
	gl_max_rectangle_texture_size_arb                     = int(0x84F8)
	gl_max_rectangle_texture_size_nv                      = int(0x84F8)
	gl_depth_stencil                                      = int(0x84F9)
	gl_depth_stencil_ext                                  = int(0x84F9)
	gl_depth_stencil_nv                                   = int(0x84F9)
	gl_depth_stencil_oes                                  = int(0x84F9)
	gl_unsigned_int_24_8                                  = int(0x84FA)
	gl_unsigned_int_24_8_ext                              = int(0x84FA)
	gl_unsigned_int_24_8_nv                               = int(0x84FA)
	gl_unsigned_int_24_8_oes                              = int(0x84FA)
	gl_max_texture_lod_bias                               = int(0x84FD)
	gl_max_texture_lod_bias_ext                           = int(0x84FD)
	gl_texture_max_anisotropy                             = int(0x84FE)
	gl_texture_max_anisotropy_ext                         = int(0x84FE)
	gl_max_texture_max_anisotropy                         = int(0x84FF)
	gl_max_texture_max_anisotropy_ext                     = int(0x84FF)
	gl_texture_filter_control                             = int(0x8500)
	gl_texture_filter_control_ext                         = int(0x8500)
	gl_texture_lod_bias                                   = int(0x8501)
	gl_texture_lod_bias_ext                               = int(0x8501)
	gl_modelview1_stack_depth_ext                         = int(0x8502)
	gl_combine4_nv                                        = int(0x8503)
	gl_max_shininess_nv                                   = int(0x8504)
	gl_max_spot_exponent_nv                               = int(0x8505)
	gl_modelview1_matrix_ext                              = int(0x8506)
	gl_incr_wrap                                          = int(0x8507)
	gl_incr_wrap_ext                                      = int(0x8507)
	gl_incr_wrap_oes                                      = int(0x8507)
	gl_decr_wrap                                          = int(0x8508)
	gl_decr_wrap_ext                                      = int(0x8508)
	gl_decr_wrap_oes                                      = int(0x8508)
	gl_vertex_weighting_ext                               = int(0x8509)
	gl_modelview1_arb                                     = int(0x850A)
	gl_modelview1_ext                                     = int(0x850A)
	gl_current_vertex_weight_ext                          = int(0x850B)
	gl_vertex_weight_array_ext                            = int(0x850C)
	gl_vertex_weight_array_size_ext                       = int(0x850D)
	gl_vertex_weight_array_type_ext                       = int(0x850E)
	gl_vertex_weight_array_stride_ext                     = int(0x850F)
	gl_vertex_weight_array_pointer_ext                    = int(0x8510)
	gl_normal_map                                         = int(0x8511)
	gl_normal_map_arb                                     = int(0x8511)
	gl_normal_map_ext                                     = int(0x8511)
	gl_normal_map_nv                                      = int(0x8511)
	gl_normal_map_oes                                     = int(0x8511)
	gl_reflection_map                                     = int(0x8512)
	gl_reflection_map_arb                                 = int(0x8512)
	gl_reflection_map_ext                                 = int(0x8512)
	gl_reflection_map_nv                                  = int(0x8512)
	gl_reflection_map_oes                                 = int(0x8512)
	gl_texture_cube_map                                   = int(0x8513)
	gl_texture_cube_map_arb                               = int(0x8513)
	gl_texture_cube_map_ext                               = int(0x8513)
	gl_texture_cube_map_oes                               = int(0x8513)
	gl_texture_binding_cube_map                           = int(0x8514)
	gl_texture_binding_cube_map_arb                       = int(0x8514)
	gl_texture_binding_cube_map_ext                       = int(0x8514)
	gl_texture_binding_cube_map_oes                       = int(0x8514)
	gl_texture_cube_map_positive_x                        = int(0x8515)
	gl_texture_cube_map_positive_x_arb                    = int(0x8515)
	gl_texture_cube_map_positive_x_ext                    = int(0x8515)
	gl_texture_cube_map_positive_x_oes                    = int(0x8515)
	gl_texture_cube_map_negative_x                        = int(0x8516)
	gl_texture_cube_map_negative_x_arb                    = int(0x8516)
	gl_texture_cube_map_negative_x_ext                    = int(0x8516)
	gl_texture_cube_map_negative_x_oes                    = int(0x8516)
	gl_texture_cube_map_positive_y                        = int(0x8517)
	gl_texture_cube_map_positive_y_arb                    = int(0x8517)
	gl_texture_cube_map_positive_y_ext                    = int(0x8517)
	gl_texture_cube_map_positive_y_oes                    = int(0x8517)
	gl_texture_cube_map_negative_y                        = int(0x8518)
	gl_texture_cube_map_negative_y_arb                    = int(0x8518)
	gl_texture_cube_map_negative_y_ext                    = int(0x8518)
	gl_texture_cube_map_negative_y_oes                    = int(0x8518)
	gl_texture_cube_map_positive_z                        = int(0x8519)
	gl_texture_cube_map_positive_z_arb                    = int(0x8519)
	gl_texture_cube_map_positive_z_ext                    = int(0x8519)
	gl_texture_cube_map_positive_z_oes                    = int(0x8519)
	gl_texture_cube_map_negative_z                        = int(0x851A)
	gl_texture_cube_map_negative_z_arb                    = int(0x851A)
	gl_texture_cube_map_negative_z_ext                    = int(0x851A)
	gl_texture_cube_map_negative_z_oes                    = int(0x851A)
	gl_proxy_texture_cube_map                             = int(0x851B)
	gl_proxy_texture_cube_map_arb                         = int(0x851B)
	gl_proxy_texture_cube_map_ext                         = int(0x851B)
	gl_max_cube_map_texture_size                          = int(0x851C)
	gl_max_cube_map_texture_size_arb                      = int(0x851C)
	gl_max_cube_map_texture_size_ext                      = int(0x851C)
	gl_max_cube_map_texture_size_oes                      = int(0x851C)
	gl_vertex_array_range_apple                           = int(0x851D)
	gl_vertex_array_range_nv                              = int(0x851D)
	gl_vertex_array_range_length_apple                    = int(0x851E)
	gl_vertex_array_range_length_nv                       = int(0x851E)
	gl_vertex_array_range_valid_nv                        = int(0x851F)
	gl_vertex_array_storage_hint_apple                    = int(0x851F)
	gl_max_vertex_array_range_element_nv                  = int(0x8520)
	gl_vertex_array_range_pointer_apple                   = int(0x8521)
	gl_vertex_array_range_pointer_nv                      = int(0x8521)
	gl_register_combiners_nv                              = int(0x8522)
	gl_variable_a_nv                                      = int(0x8523)
	gl_variable_b_nv                                      = int(0x8524)
	gl_variable_c_nv                                      = int(0x8525)
	gl_variable_d_nv                                      = int(0x8526)
	gl_variable_e_nv                                      = int(0x8527)
	gl_variable_f_nv                                      = int(0x8528)
	gl_variable_g_nv                                      = int(0x8529)
	gl_constant_color0_nv                                 = int(0x852A)
	gl_constant_color1_nv                                 = int(0x852B)
	gl_primary_color_nv                                   = int(0x852C)
	gl_secondary_color_nv                                 = int(0x852D)
	gl_spare0_nv                                          = int(0x852E)
	gl_spare1_nv                                          = int(0x852F)
	gl_discard_nv                                         = int(0x8530)
	gl_e_times_f_nv                                       = int(0x8531)
	gl_spare0_plus_secondary_color_nv                     = int(0x8532)
	gl_vertex_array_range_without_flush_nv                = int(0x8533)
	gl_multisample_filter_hint_nv                         = int(0x8534)
	gl_per_stage_constants_nv                             = int(0x8535)
	gl_unsigned_identity_nv                               = int(0x8536)
	gl_unsigned_invert_nv                                 = int(0x8537)
	gl_expand_normal_nv                                   = int(0x8538)
	gl_expand_negate_nv                                   = int(0x8539)
	gl_half_bias_normal_nv                                = int(0x853A)
	gl_half_bias_negate_nv                                = int(0x853B)
	gl_signed_identity_nv                                 = int(0x853C)
	gl_signed_negate_nv                                   = int(0x853D)
	gl_scale_by_two_nv                                    = int(0x853E)
	gl_scale_by_four_nv                                   = int(0x853F)
	gl_scale_by_one_half_nv                               = int(0x8540)
	gl_bias_by_negative_one_half_nv                       = int(0x8541)
	gl_combiner_input_nv                                  = int(0x8542)
	gl_combiner_mapping_nv                                = int(0x8543)
	gl_combiner_component_usage_nv                        = int(0x8544)
	gl_combiner_ab_dot_product_nv                         = int(0x8545)
	gl_combiner_cd_dot_product_nv                         = int(0x8546)
	gl_combiner_mux_sum_nv                                = int(0x8547)
	gl_combiner_scale_nv                                  = int(0x8548)
	gl_combiner_bias_nv                                   = int(0x8549)
	gl_combiner_ab_output_nv                              = int(0x854A)
	gl_combiner_cd_output_nv                              = int(0x854B)
	gl_combiner_sum_output_nv                             = int(0x854C)
	gl_max_general_combiners_nv                           = int(0x854D)
	gl_num_general_combiners_nv                           = int(0x854E)
	gl_color_sum_clamp_nv                                 = int(0x854F)
	gl_combiner0_nv                                       = int(0x8550)
	gl_combiner1_nv                                       = int(0x8551)
	gl_combiner2_nv                                       = int(0x8552)
	gl_combiner3_nv                                       = int(0x8553)
	gl_combiner4_nv                                       = int(0x8554)
	gl_combiner5_nv                                       = int(0x8555)
	gl_combiner6_nv                                       = int(0x8556)
	gl_combiner7_nv                                       = int(0x8557)
	gl_primitive_restart_nv                               = int(0x8558)
	gl_primitive_restart_index_nv                         = int(0x8559)
	gl_fog_distance_mode_nv                               = int(0x855A)
	gl_eye_radial_nv                                      = int(0x855B)
	gl_eye_plane_absolute_nv                              = int(0x855C)
	gl_emboss_light_nv                                    = int(0x855D)
	gl_emboss_constant_nv                                 = int(0x855E)
	gl_emboss_map_nv                                      = int(0x855F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8560" end="0x856F" vendor="ZiiLabs" |>
pub const (
	gl_red_min_clamp_ingr   = int(0x8560)
	gl_green_min_clamp_ingr = int(0x8561)
	gl_blue_min_clamp_ingr  = int(0x8562)
	gl_alpha_min_clamp_ingr = int(0x8563)
	gl_red_max_clamp_ingr   = int(0x8564)
	gl_green_max_clamp_ingr = int(0x8565)
	gl_blue_max_clamp_ingr  = int(0x8566)
	gl_alpha_max_clamp_ingr = int(0x8567)
	gl_interlace_read_ingr  = int(0x8568)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8570" end="0x859F" group="TextureEnvParameter" vendor="AMD/NV" |>
pub const (
	gl_combine            = int(0x8570)
	gl_combine_arb        = int(0x8570)
	gl_combine_ext        = int(0x8570)
	gl_combine_rgb        = int(0x8571)
	gl_combine_rgb_arb    = int(0x8571)
	gl_combine_rgb_ext    = int(0x8571)
	gl_combine_alpha      = int(0x8572)
	gl_combine_alpha_arb  = int(0x8572)
	gl_combine_alpha_ext  = int(0x8572)
	gl_rgb_scale          = int(0x8573)
	gl_rgb_scale_arb      = int(0x8573)
	gl_rgb_scale_ext      = int(0x8573)
	gl_add_signed         = int(0x8574)
	gl_add_signed_arb     = int(0x8574)
	gl_add_signed_ext     = int(0x8574)
	gl_interpolate        = int(0x8575)
	gl_interpolate_arb    = int(0x8575)
	gl_interpolate_ext    = int(0x8575)
	gl_constant           = int(0x8576)
	gl_constant_arb       = int(0x8576)
	gl_constant_ext       = int(0x8576)
	gl_constant_nv        = int(0x8576)
	gl_primary_color      = int(0x8577)
	gl_primary_color_arb  = int(0x8577)
	gl_primary_color_ext  = int(0x8577)
	gl_previous           = int(0x8578)
	gl_previous_arb       = int(0x8578)
	gl_previous_ext       = int(0x8578)
	gl_source0_rgb        = int(0x8580)
	gl_source0_rgb_arb    = int(0x8580)
	gl_source0_rgb_ext    = int(0x8580)
	gl_src0_rgb           = int(0x8580)
	gl_source1_rgb        = int(0x8581)
	gl_source1_rgb_arb    = int(0x8581)
	gl_source1_rgb_ext    = int(0x8581)
	gl_src1_rgb           = int(0x8581)
	gl_source2_rgb        = int(0x8582)
	gl_source2_rgb_arb    = int(0x8582)
	gl_source2_rgb_ext    = int(0x8582)
	gl_src2_rgb           = int(0x8582)
	gl_source3_rgb_nv     = int(0x8583)
	gl_source0_alpha      = int(0x8588)
	gl_source0_alpha_arb  = int(0x8588)
	gl_source0_alpha_ext  = int(0x8588)
	gl_src0_alpha         = int(0x8588)
	gl_source1_alpha      = int(0x8589)
	gl_source1_alpha_arb  = int(0x8589)
	gl_source1_alpha_ext  = int(0x8589)
	gl_src1_alpha         = int(0x8589)
	gl_src1_alpha_ext     = int(0x8589)
	gl_source2_alpha      = int(0x858A)
	gl_source2_alpha_arb  = int(0x858A)
	gl_source2_alpha_ext  = int(0x858A)
	gl_src2_alpha         = int(0x858A)
	gl_source3_alpha_nv   = int(0x858B)
	gl_operand0_rgb       = int(0x8590)
	gl_operand0_rgb_arb   = int(0x8590)
	gl_operand0_rgb_ext   = int(0x8590)
	gl_operand1_rgb       = int(0x8591)
	gl_operand1_rgb_arb   = int(0x8591)
	gl_operand1_rgb_ext   = int(0x8591)
	gl_operand2_rgb       = int(0x8592)
	gl_operand2_rgb_arb   = int(0x8592)
	gl_operand2_rgb_ext   = int(0x8592)
	gl_operand3_rgb_nv    = int(0x8593)
	gl_operand0_alpha     = int(0x8598)
	gl_operand0_alpha_arb = int(0x8598)
	gl_operand0_alpha_ext = int(0x8598)
	gl_operand1_alpha     = int(0x8599)
	gl_operand1_alpha_arb = int(0x8599)
	gl_operand1_alpha_ext = int(0x8599)
	gl_operand2_alpha     = int(0x859A)
	gl_operand2_alpha_arb = int(0x859A)
	gl_operand2_alpha_ext = int(0x859A)
	gl_operand3_alpha_nv  = int(0x859B)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x85A0" end="0x85AF" vendor="SGI" |>
pub const (
	gl_pack_subsample_rate_sgix   = int(0x85A0)
	gl_unpack_subsample_rate_sgix = int(0x85A1)
	gl_pixel_subsample_4444_sgix  = int(0x85A2)
	gl_pixel_subsample_2424_sgix  = int(0x85A3)
	gl_pixel_subsample_4242_sgix  = int(0x85A4)
	gl_perturb_ext                = int(0x85AE)
	gl_texture_normal_ext         = int(0x85AF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x85B0" end="0x85BF" vendor="APPLE" |>
pub const (
	gl_light_model_specular_vector_apple = int(0x85B0)
	gl_transform_hint_apple              = int(0x85B1)
	gl_unpack_client_storage_apple       = int(0x85B2)
	gl_buffer_object_apple               = int(0x85B3)
	gl_storage_client_apple              = int(0x85B4)
	gl_vertex_array_binding              = int(0x85B5)
	gl_vertex_array_binding_apple        = int(0x85B5)
	gl_vertex_array_binding_oes          = int(0x85B5)
	gl_texture_range_length_apple        = int(0x85B7)
	gl_texture_range_pointer_apple       = int(0x85B8)
	gl_ycbcr_422_apple                   = int(0x85B9)
	gl_unsigned_short_8_8_apple          = int(0x85BA)
	gl_unsigned_short_8_8_mesa           = int(0x85BA)
	gl_unsigned_short_8_8_rev_apple      = int(0x85BB)
	gl_unsigned_short_8_8_rev_mesa       = int(0x85BB)
	gl_texture_storage_hint_apple        = int(0x85BC)
	gl_storage_private_apple             = int(0x85BD)
	gl_storage_cached_apple              = int(0x85BE)
	gl_storage_shared_apple              = int(0x85BF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x85C0" end="0x85CF" vendor="SUN" |>
pub const (
	gl_replacement_code_array_sun         = int(0x85C0)
	gl_replacement_code_array_type_sun    = int(0x85C1)
	gl_replacement_code_array_stride_sun  = int(0x85C2)
	gl_replacement_code_array_pointer_sun = int(0x85C3)
	gl_r1ui_v3f_sun                       = int(0x85C4)
	gl_r1ui_c4ub_v3f_sun                  = int(0x85C5)
	gl_r1ui_c3f_v3f_sun                   = int(0x85C6)
	gl_r1ui_n3f_v3f_sun                   = int(0x85C7)
	gl_r1ui_c4f_n3f_v3f_sun               = int(0x85C8)
	gl_r1ui_t2f_v3f_sun                   = int(0x85C9)
	gl_r1ui_t2f_n3f_v3f_sun               = int(0x85CA)
	gl_r1ui_t2f_c4f_n3f_v3f_sun           = int(0x85CB)
	gl_slice_accum_sun                    = int(0x85CC)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8600" end="0x861F" vendor="SUN" |>
pub const (
	gl_quad_mesh_sun     = int(0x8614)
	gl_triangle_mesh_sun = int(0x8615)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8620" end="0x867F" vendor="NV" |>
pub const (
	gl_vertex_program_arb                 = int(0x8620)
	gl_vertex_program_nv                  = int(0x8620)
	gl_vertex_state_program_nv            = int(0x8621)
	gl_vertex_attrib_array_enabled        = int(0x8622)
	gl_vertex_attrib_array_enabled_arb    = int(0x8622)
	gl_attrib_array_size_nv               = int(0x8623)
	gl_vertex_attrib_array_size           = int(0x8623)
	gl_vertex_attrib_array_size_arb       = int(0x8623)
	gl_attrib_array_stride_nv             = int(0x8624)
	gl_vertex_attrib_array_stride         = int(0x8624)
	gl_vertex_attrib_array_stride_arb     = int(0x8624)
	gl_attrib_array_type_nv               = int(0x8625)
	gl_vertex_attrib_array_type           = int(0x8625)
	gl_vertex_attrib_array_type_arb       = int(0x8625)
	gl_current_attrib_nv                  = int(0x8626)
	gl_current_vertex_attrib              = int(0x8626)
	gl_current_vertex_attrib_arb          = int(0x8626)
	gl_program_length_arb                 = int(0x8627)
	gl_program_length_nv                  = int(0x8627)
	gl_program_string_arb                 = int(0x8628)
	gl_program_string_nv                  = int(0x8628)
	gl_modelview_projection_nv            = int(0x8629)
	gl_identity_nv                        = int(0x862A)
	gl_inverse_nv                         = int(0x862B)
	gl_transpose_nv                       = int(0x862C)
	gl_inverse_transpose_nv               = int(0x862D)
	gl_max_program_matrix_stack_depth_arb = int(0x862E)
	gl_max_track_matrix_stack_depth_nv    = int(0x862E)
	gl_max_program_matrices_arb           = int(0x862F)
	gl_max_track_matrices_nv              = int(0x862F)
	gl_matrix0_nv                         = int(0x8630)
	gl_matrix1_nv                         = int(0x8631)
	gl_matrix2_nv                         = int(0x8632)
	gl_matrix3_nv                         = int(0x8633)
	gl_matrix4_nv                         = int(0x8634)
	gl_matrix5_nv                         = int(0x8635)
	gl_matrix6_nv                         = int(0x8636)
	gl_matrix7_nv                         = int(0x8637)
	gl_current_matrix_stack_depth_arb     = int(0x8640)
	gl_current_matrix_stack_depth_nv      = int(0x8640)
	gl_current_matrix_arb                 = int(0x8641)
	gl_current_matrix_nv                  = int(0x8641)
	gl_vertex_program_point_size          = int(0x8642)
	gl_vertex_program_point_size_arb      = int(0x8642)
	gl_vertex_program_point_size_nv       = int(0x8642)
	gl_program_point_size                 = int(0x8642)
	gl_program_point_size_arb             = int(0x8642)
	gl_program_point_size_ext             = int(0x8642)
	gl_vertex_program_two_side            = int(0x8643)
	gl_vertex_program_two_side_arb        = int(0x8643)
	gl_vertex_program_two_side_nv         = int(0x8643)
	gl_program_parameter_nv               = int(0x8644)
	gl_attrib_array_pointer_nv            = int(0x8645)
	gl_vertex_attrib_array_pointer        = int(0x8645)
	gl_vertex_attrib_array_pointer_arb    = int(0x8645)
	gl_program_target_nv                  = int(0x8646)
	gl_program_resident_nv                = int(0x8647)
	gl_track_matrix_nv                    = int(0x8648)
	gl_track_matrix_transform_nv          = int(0x8649)
	gl_vertex_program_binding_nv          = int(0x864A)
	gl_program_error_position_arb         = int(0x864B)
	gl_program_error_position_nv          = int(0x864B)
	gl_offset_texture_rectangle_nv        = int(0x864C)
	gl_offset_texture_rectangle_scale_nv  = int(0x864D)
	gl_dot_product_texture_rectangle_nv   = int(0x864E)
	gl_depth_clamp                        = int(0x864F)
	gl_depth_clamp_nv                     = int(0x864F)
	gl_depth_clamp_ext                    = int(0x864F)
	gl_vertex_attrib_array0_nv            = int(0x8650)
	gl_vertex_attrib_array1_nv            = int(0x8651)
	gl_vertex_attrib_array2_nv            = int(0x8652)
	gl_vertex_attrib_array3_nv            = int(0x8653)
	gl_vertex_attrib_array4_nv            = int(0x8654)
	gl_vertex_attrib_array5_nv            = int(0x8655)
	gl_vertex_attrib_array6_nv            = int(0x8656)
	gl_vertex_attrib_array7_nv            = int(0x8657)
	gl_vertex_attrib_array8_nv            = int(0x8658)
	gl_vertex_attrib_array9_nv            = int(0x8659)
	gl_vertex_attrib_array10_nv           = int(0x865A)
	gl_vertex_attrib_array11_nv           = int(0x865B)
	gl_vertex_attrib_array12_nv           = int(0x865C)
	gl_vertex_attrib_array13_nv           = int(0x865D)
	gl_vertex_attrib_array14_nv           = int(0x865E)
	gl_vertex_attrib_array15_nv           = int(0x865F)
	gl_map1_vertex_attrib0_4_nv           = int(0x8660)
	gl_map1_vertex_attrib1_4_nv           = int(0x8661)
	gl_map1_vertex_attrib2_4_nv           = int(0x8662)
	gl_map1_vertex_attrib3_4_nv           = int(0x8663)
	gl_map1_vertex_attrib4_4_nv           = int(0x8664)
	gl_map1_vertex_attrib5_4_nv           = int(0x8665)
	gl_map1_vertex_attrib6_4_nv           = int(0x8666)
	gl_map1_vertex_attrib7_4_nv           = int(0x8667)
	gl_map1_vertex_attrib8_4_nv           = int(0x8668)
	gl_map1_vertex_attrib9_4_nv           = int(0x8669)
	gl_map1_vertex_attrib10_4_nv          = int(0x866A)
	gl_map1_vertex_attrib11_4_nv          = int(0x866B)
	gl_map1_vertex_attrib12_4_nv          = int(0x866C)
	gl_map1_vertex_attrib13_4_nv          = int(0x866D)
	gl_map1_vertex_attrib14_4_nv          = int(0x866E)
	gl_map1_vertex_attrib15_4_nv          = int(0x866F)
	gl_map2_vertex_attrib0_4_nv           = int(0x8670)
	gl_map2_vertex_attrib1_4_nv           = int(0x8671)
	gl_map2_vertex_attrib2_4_nv           = int(0x8672)
	gl_map2_vertex_attrib3_4_nv           = int(0x8673)
	gl_map2_vertex_attrib4_4_nv           = int(0x8674)
	gl_map2_vertex_attrib5_4_nv           = int(0x8675)
	gl_map2_vertex_attrib6_4_nv           = int(0x8676)
	gl_map2_vertex_attrib7_4_nv           = int(0x8677)
	gl_program_binding_arb                = int(0x8677)
	gl_map2_vertex_attrib8_4_nv           = int(0x8678)
	gl_map2_vertex_attrib9_4_nv           = int(0x8679)
	gl_map2_vertex_attrib10_4_nv          = int(0x867A)
	gl_map2_vertex_attrib11_4_nv          = int(0x867B)
	gl_map2_vertex_attrib12_4_nv          = int(0x867C)
	gl_map2_vertex_attrib13_4_nv          = int(0x867D)
	gl_map2_vertex_attrib14_4_nv          = int(0x867E)
	gl_map2_vertex_attrib15_4_nv          = int(0x867F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x86A0" end="0x86AF" vendor="ARB" |>
pub const (
	gl_texture_compressed_image_size      = int(0x86A0)
	gl_texture_compressed_image_size_arb  = int(0x86A0)
	gl_texture_compressed                 = int(0x86A1)
	gl_texture_compressed_arb             = int(0x86A1)
	gl_num_compressed_texture_formats     = int(0x86A2)
	gl_num_compressed_texture_formats_arb = int(0x86A2)
	gl_compressed_texture_formats         = int(0x86A3)
	gl_compressed_texture_formats_arb     = int(0x86A3)
	gl_max_vertex_units_arb               = int(0x86A4)
	gl_max_vertex_units_oes               = int(0x86A4)
	gl_active_vertex_units_arb            = int(0x86A5)
	gl_weight_sum_unity_arb               = int(0x86A6)
	gl_vertex_blend_arb                   = int(0x86A7)
	gl_current_weight_arb                 = int(0x86A8)
	gl_weight_array_type_arb              = int(0x86A9)
	gl_weight_array_type_oes              = int(0x86A9)
	gl_weight_array_stride_arb            = int(0x86AA)
	gl_weight_array_stride_oes            = int(0x86AA)
	gl_weight_array_size_arb              = int(0x86AB)
	gl_weight_array_size_oes              = int(0x86AB)
	gl_weight_array_pointer_arb           = int(0x86AC)
	gl_weight_array_pointer_oes           = int(0x86AC)
	gl_weight_array_arb                   = int(0x86AD)
	gl_weight_array_oes                   = int(0x86AD)
	gl_dot3_rgb                           = int(0x86AE)
	gl_dot3_rgb_arb                       = int(0x86AE)
	gl_dot3_rgba                          = int(0x86AF)
	gl_dot3_rgba_arb                      = int(0x86AF)
	gl_dot3_rgba_img                      = int(0x86AF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x86B0" end="0x86BF" vendor="3DFX" |>
pub const (
	gl_compressed_rgb_fxt1_3dfx  = int(0x86B0)
	gl_compressed_rgba_fxt1_3dfx = int(0x86B1)
	gl_multisample_3dfx          = int(0x86B2)
	gl_sample_buffers_3dfx       = int(0x86B3)
	gl_samples_3dfx              = int(0x86B4)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x86C0" end="0x871F" vendor="NV" |>
pub const (
	gl_eval_2d_nv                                = int(0x86C0)
	gl_eval_triangular_2d_nv                     = int(0x86C1)
	gl_map_tessellation_nv                       = int(0x86C2)
	gl_map_attrib_u_order_nv                     = int(0x86C3)
	gl_map_attrib_v_order_nv                     = int(0x86C4)
	gl_eval_fractional_tessellation_nv           = int(0x86C5)
	gl_eval_vertex_attrib0_nv                    = int(0x86C6)
	gl_eval_vertex_attrib1_nv                    = int(0x86C7)
	gl_eval_vertex_attrib2_nv                    = int(0x86C8)
	gl_eval_vertex_attrib3_nv                    = int(0x86C9)
	gl_eval_vertex_attrib4_nv                    = int(0x86CA)
	gl_eval_vertex_attrib5_nv                    = int(0x86CB)
	gl_eval_vertex_attrib6_nv                    = int(0x86CC)
	gl_eval_vertex_attrib7_nv                    = int(0x86CD)
	gl_eval_vertex_attrib8_nv                    = int(0x86CE)
	gl_eval_vertex_attrib9_nv                    = int(0x86CF)
	gl_eval_vertex_attrib10_nv                   = int(0x86D0)
	gl_eval_vertex_attrib11_nv                   = int(0x86D1)
	gl_eval_vertex_attrib12_nv                   = int(0x86D2)
	gl_eval_vertex_attrib13_nv                   = int(0x86D3)
	gl_eval_vertex_attrib14_nv                   = int(0x86D4)
	gl_eval_vertex_attrib15_nv                   = int(0x86D5)
	gl_max_map_tessellation_nv                   = int(0x86D6)
	gl_max_rational_eval_order_nv                = int(0x86D7)
	gl_max_program_patch_attribs_nv              = int(0x86D8)
	gl_rgba_unsigned_dot_product_mapping_nv      = int(0x86D9)
	gl_unsigned_int_s8_s8_8_8_nv                 = int(0x86DA)
	gl_unsigned_int_8_8_s8_s8_rev_nv             = int(0x86DB)
	gl_dsdt_mag_intensity_nv                     = int(0x86DC)
	gl_shader_consistent_nv                      = int(0x86DD)
	gl_texture_shader_nv                         = int(0x86DE)
	gl_shader_operation_nv                       = int(0x86DF)
	gl_cull_modes_nv                             = int(0x86E0)
	gl_offset_texture_matrix_nv                  = int(0x86E1)
	gl_offset_texture_2d_matrix_nv               = int(0x86E1)
	gl_offset_texture_scale_nv                   = int(0x86E2)
	gl_offset_texture_2d_scale_nv                = int(0x86E2)
	gl_offset_texture_bias_nv                    = int(0x86E3)
	gl_offset_texture_2d_bias_nv                 = int(0x86E3)
	gl_previous_texture_input_nv                 = int(0x86E4)
	gl_const_eye_nv                              = int(0x86E5)
	gl_pass_through_nv                           = int(0x86E6)
	gl_cull_fragment_nv                          = int(0x86E7)
	gl_offset_texture_2d_nv                      = int(0x86E8)
	gl_dependent_ar_texture_2d_nv                = int(0x86E9)
	gl_dependent_gb_texture_2d_nv                = int(0x86EA)
	gl_surface_state_nv                          = int(0x86EB)
	gl_dot_product_nv                            = int(0x86EC)
	gl_dot_product_depth_replace_nv              = int(0x86ED)
	gl_dot_product_texture_2d_nv                 = int(0x86EE)
	gl_dot_product_texture_3d_nv                 = int(0x86EF)
	gl_dot_product_texture_cube_map_nv           = int(0x86F0)
	gl_dot_product_diffuse_cube_map_nv           = int(0x86F1)
	gl_dot_product_reflect_cube_map_nv           = int(0x86F2)
	gl_dot_product_const_eye_reflect_cube_map_nv = int(0x86F3)
	gl_hilo_nv                                   = int(0x86F4)
	gl_dsdt_nv                                   = int(0x86F5)
	gl_dsdt_mag_nv                               = int(0x86F6)
	gl_dsdt_mag_vib_nv                           = int(0x86F7)
	gl_hilo16_nv                                 = int(0x86F8)
	gl_signed_hilo_nv                            = int(0x86F9)
	gl_signed_hilo16_nv                          = int(0x86FA)
	gl_signed_rgba_nv                            = int(0x86FB)
	gl_signed_rgba8_nv                           = int(0x86FC)
	gl_surface_registered_nv                     = int(0x86FD)
	gl_signed_rgb_nv                             = int(0x86FE)
	gl_signed_rgb8_nv                            = int(0x86FF)
	gl_surface_mapped_nv                         = int(0x8700)
	gl_signed_luminance_nv                       = int(0x8701)
	gl_signed_luminance8_nv                      = int(0x8702)
	gl_signed_luminance_alpha_nv                 = int(0x8703)
	gl_signed_luminance8_alpha8_nv               = int(0x8704)
	gl_signed_alpha_nv                           = int(0x8705)
	gl_signed_alpha8_nv                          = int(0x8706)
	gl_signed_intensity_nv                       = int(0x8707)
	gl_signed_intensity8_nv                      = int(0x8708)
	gl_dsdt8_nv                                  = int(0x8709)
	gl_dsdt8_mag8_nv                             = int(0x870A)
	gl_dsdt8_mag8_intensity8_nv                  = int(0x870B)
	gl_signed_rgb_unsigned_alpha_nv              = int(0x870C)
	gl_signed_rgb8_unsigned_alpha8_nv            = int(0x870D)
	gl_hi_scale_nv                               = int(0x870E)
	gl_lo_scale_nv                               = int(0x870F)
	gl_ds_scale_nv                               = int(0x8710)
	gl_dt_scale_nv                               = int(0x8711)
	gl_magnitude_scale_nv                        = int(0x8712)
	gl_vibrance_scale_nv                         = int(0x8713)
	gl_hi_bias_nv                                = int(0x8714)
	gl_lo_bias_nv                                = int(0x8715)
	gl_ds_bias_nv                                = int(0x8716)
	gl_dt_bias_nv                                = int(0x8717)
	gl_magnitude_bias_nv                         = int(0x8718)
	gl_vibrance_bias_nv                          = int(0x8719)
	gl_texture_border_values_nv                  = int(0x871A)
	gl_texture_hi_size_nv                        = int(0x871B)
	gl_texture_lo_size_nv                        = int(0x871C)
	gl_texture_ds_size_nv                        = int(0x871D)
	gl_texture_dt_size_nv                        = int(0x871E)
	gl_texture_mag_size_nv                       = int(0x871F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8720" end="0x873F" vendor="ARB" |>
pub const (
	gl_modelview2_arb  = int(0x8722)
	gl_modelview3_arb  = int(0x8723)
	gl_modelview4_arb  = int(0x8724)
	gl_modelview5_arb  = int(0x8725)
	gl_modelview6_arb  = int(0x8726)
	gl_modelview7_arb  = int(0x8727)
	gl_modelview8_arb  = int(0x8728)
	gl_modelview9_arb  = int(0x8729)
	gl_modelview10_arb = int(0x872A)
	gl_modelview11_arb = int(0x872B)
	gl_modelview12_arb = int(0x872C)
	gl_modelview13_arb = int(0x872D)
	gl_modelview14_arb = int(0x872E)
	gl_modelview15_arb = int(0x872F)
	gl_modelview16_arb = int(0x8730)
	gl_modelview17_arb = int(0x8731)
	gl_modelview18_arb = int(0x8732)
	gl_modelview19_arb = int(0x8733)
	gl_modelview20_arb = int(0x8734)
	gl_modelview21_arb = int(0x8735)
	gl_modelview22_arb = int(0x8736)
	gl_modelview23_arb = int(0x8737)
	gl_modelview24_arb = int(0x8738)
	gl_modelview25_arb = int(0x8739)
	gl_modelview26_arb = int(0x873A)
	gl_modelview27_arb = int(0x873B)
	gl_modelview28_arb = int(0x873C)
	gl_modelview29_arb = int(0x873D)
	gl_modelview30_arb = int(0x873E)
	gl_modelview31_arb = int(0x873F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8740" end="0x874F" vendor="AMD" |>
pub const (
	gl_dot3_rgb_ext                   = int(0x8740)
	gl_z400_binary_amd                = int(0x8740)
	gl_dot3_rgba_ext                  = int(0x8741)
	gl_program_binary_length_oes      = int(0x8741)
	gl_program_binary_length          = int(0x8741)
	gl_mirror_clamp_ati               = int(0x8742)
	gl_mirror_clamp_ext               = int(0x8742)
	gl_mirror_clamp_to_edge           = int(0x8743)
	gl_mirror_clamp_to_edge_ati       = int(0x8743)
	gl_mirror_clamp_to_edge_ext       = int(0x8743)
	gl_modulate_add_ati               = int(0x8744)
	gl_modulate_signed_add_ati        = int(0x8745)
	gl_modulate_subtract_ati          = int(0x8746)
	gl_set_amd                        = int(0x874A)
	gl_replace_value_amd              = int(0x874B)
	gl_stencil_op_value_amd           = int(0x874C)
	gl_stencil_back_op_value_amd      = int(0x874D)
	gl_vertex_attrib_array_long       = int(0x874E)
	gl_occlusion_query_event_mask_amd = int(0x874F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8750" end="0x875F" vendor="MESA" |>
pub const (
	gl_depth_stencil_mesa             = int(0x8750)
	gl_unsigned_int_24_8_mesa         = int(0x8751)
	gl_unsigned_int_8_24_rev_mesa     = int(0x8752)
	gl_unsigned_short_15_1_mesa       = int(0x8753)
	gl_unsigned_short_1_15_rev_mesa   = int(0x8754)
	gl_trace_mask_mesa                = int(0x8755)
	gl_trace_name_mesa                = int(0x8756)
	gl_ycbcr_mesa                     = int(0x8757)
	gl_pack_invert_mesa               = int(0x8758)
	gl_debug_object_mesa              = int(0x8759)
	gl_texture_1d_stack_mesax         = int(0x8759)
	gl_debug_print_mesa               = int(0x875A)
	gl_texture_2d_stack_mesax         = int(0x875A)
	gl_debug_assert_mesa              = int(0x875B)
	gl_proxy_texture_1d_stack_mesax   = int(0x875B)
	gl_proxy_texture_2d_stack_mesax   = int(0x875C)
	gl_texture_1d_stack_binding_mesax = int(0x875D)
	gl_texture_2d_stack_binding_mesax = int(0x875E)
	gl_program_binary_format_mesa     = int(0x875F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8760" end="0x883F" vendor="AMD" |>
pub const (
	gl_static_ati                                      = int(0x8760)
	gl_dynamic_ati                                     = int(0x8761)
	gl_preserve_ati                                    = int(0x8762)
	gl_discard_ati                                     = int(0x8763)
	gl_buffer_size                                     = int(0x8764)
	gl_buffer_size_arb                                 = int(0x8764)
	gl_object_buffer_size_ati                          = int(0x8764)
	gl_buffer_usage                                    = int(0x8765)
	gl_buffer_usage_arb                                = int(0x8765)
	gl_object_buffer_usage_ati                         = int(0x8765)
	gl_array_object_buffer_ati                         = int(0x8766)
	gl_array_object_offset_ati                         = int(0x8767)
	gl_element_array_ati                               = int(0x8768)
	gl_element_array_type_ati                          = int(0x8769)
	gl_element_array_pointer_ati                       = int(0x876A)
	gl_max_vertex_streams_ati                          = int(0x876B)
	gl_vertex_stream0_ati                              = int(0x876C)
	gl_vertex_stream1_ati                              = int(0x876D)
	gl_vertex_stream2_ati                              = int(0x876E)
	gl_vertex_stream3_ati                              = int(0x876F)
	gl_vertex_stream4_ati                              = int(0x8770)
	gl_vertex_stream5_ati                              = int(0x8771)
	gl_vertex_stream6_ati                              = int(0x8772)
	gl_vertex_stream7_ati                              = int(0x8773)
	gl_vertex_source_ati                               = int(0x8774)
	gl_bump_rot_matrix_ati                             = int(0x8775)
	gl_bump_rot_matrix_size_ati                        = int(0x8776)
	gl_bump_num_tex_units_ati                          = int(0x8777)
	gl_bump_tex_units_ati                              = int(0x8778)
	gl_dudv_ati                                        = int(0x8779)
	gl_du8dv8_ati                                      = int(0x877A)
	gl_bump_envmap_ati                                 = int(0x877B)
	gl_bump_target_ati                                 = int(0x877C)
	gl_vertex_shader_ext                               = int(0x8780)
	gl_vertex_shader_binding_ext                       = int(0x8781)
	gl_op_index_ext                                    = int(0x8782)
	gl_op_negate_ext                                   = int(0x8783)
	gl_op_dot3_ext                                     = int(0x8784)
	gl_op_dot4_ext                                     = int(0x8785)
	gl_op_mul_ext                                      = int(0x8786)
	gl_op_add_ext                                      = int(0x8787)
	gl_op_madd_ext                                     = int(0x8788)
	gl_op_frac_ext                                     = int(0x8789)
	gl_op_max_ext                                      = int(0x878A)
	gl_op_min_ext                                      = int(0x878B)
	gl_op_set_ge_ext                                   = int(0x878C)
	gl_op_set_lt_ext                                   = int(0x878D)
	gl_op_clamp_ext                                    = int(0x878E)
	gl_op_floor_ext                                    = int(0x878F)
	gl_op_round_ext                                    = int(0x8790)
	gl_op_exp_base_2_ext                               = int(0x8791)
	gl_op_log_base_2_ext                               = int(0x8792)
	gl_op_power_ext                                    = int(0x8793)
	gl_op_recip_ext                                    = int(0x8794)
	gl_op_recip_sqrt_ext                               = int(0x8795)
	gl_op_sub_ext                                      = int(0x8796)
	gl_op_cross_product_ext                            = int(0x8797)
	gl_op_multiply_matrix_ext                          = int(0x8798)
	gl_op_mov_ext                                      = int(0x8799)
	gl_output_vertex_ext                               = int(0x879A)
	gl_output_color0_ext                               = int(0x879B)
	gl_output_color1_ext                               = int(0x879C)
	gl_output_texture_coord0_ext                       = int(0x879D)
	gl_output_texture_coord1_ext                       = int(0x879E)
	gl_output_texture_coord2_ext                       = int(0x879F)
	gl_output_texture_coord3_ext                       = int(0x87A0)
	gl_output_texture_coord4_ext                       = int(0x87A1)
	gl_output_texture_coord5_ext                       = int(0x87A2)
	gl_output_texture_coord6_ext                       = int(0x87A3)
	gl_output_texture_coord7_ext                       = int(0x87A4)
	gl_output_texture_coord8_ext                       = int(0x87A5)
	gl_output_texture_coord9_ext                       = int(0x87A6)
	gl_output_texture_coord10_ext                      = int(0x87A7)
	gl_output_texture_coord11_ext                      = int(0x87A8)
	gl_output_texture_coord12_ext                      = int(0x87A9)
	gl_output_texture_coord13_ext                      = int(0x87AA)
	gl_output_texture_coord14_ext                      = int(0x87AB)
	gl_output_texture_coord15_ext                      = int(0x87AC)
	gl_output_texture_coord16_ext                      = int(0x87AD)
	gl_output_texture_coord17_ext                      = int(0x87AE)
	gl_output_texture_coord18_ext                      = int(0x87AF)
	gl_output_texture_coord19_ext                      = int(0x87B0)
	gl_output_texture_coord20_ext                      = int(0x87B1)
	gl_output_texture_coord21_ext                      = int(0x87B2)
	gl_output_texture_coord22_ext                      = int(0x87B3)
	gl_output_texture_coord23_ext                      = int(0x87B4)
	gl_output_texture_coord24_ext                      = int(0x87B5)
	gl_output_texture_coord25_ext                      = int(0x87B6)
	gl_output_texture_coord26_ext                      = int(0x87B7)
	gl_output_texture_coord27_ext                      = int(0x87B8)
	gl_output_texture_coord28_ext                      = int(0x87B9)
	gl_output_texture_coord29_ext                      = int(0x87BA)
	gl_output_texture_coord30_ext                      = int(0x87BB)
	gl_output_texture_coord31_ext                      = int(0x87BC)
	gl_output_fog_ext                                  = int(0x87BD)
	gl_scalar_ext                                      = int(0x87BE)
	gl_vector_ext                                      = int(0x87BF)
	gl_matrix_ext                                      = int(0x87C0)
	gl_variant_ext                                     = int(0x87C1)
	gl_invariant_ext                                   = int(0x87C2)
	gl_local_constant_ext                              = int(0x87C3)
	gl_local_ext                                       = int(0x87C4)
	gl_max_vertex_shader_instructions_ext              = int(0x87C5)
	gl_max_vertex_shader_variants_ext                  = int(0x87C6)
	gl_max_vertex_shader_invariants_ext                = int(0x87C7)
	gl_max_vertex_shader_local_constants_ext           = int(0x87C8)
	gl_max_vertex_shader_locals_ext                    = int(0x87C9)
	gl_max_optimized_vertex_shader_instructions_ext    = int(0x87CA)
	gl_max_optimized_vertex_shader_variants_ext        = int(0x87CB)
	gl_max_optimized_vertex_shader_local_constants_ext = int(0x87CC)
	gl_max_optimized_vertex_shader_invariants_ext      = int(0x87CD)
	gl_max_optimized_vertex_shader_locals_ext          = int(0x87CE)
	gl_vertex_shader_instructions_ext                  = int(0x87CF)
	gl_vertex_shader_variants_ext                      = int(0x87D0)
	gl_vertex_shader_invariants_ext                    = int(0x87D1)
	gl_vertex_shader_local_constants_ext               = int(0x87D2)
	gl_vertex_shader_locals_ext                        = int(0x87D3)
	gl_vertex_shader_optimized_ext                     = int(0x87D4)
	gl_x_ext                                           = int(0x87D5)
	gl_y_ext                                           = int(0x87D6)
	gl_z_ext                                           = int(0x87D7)
	gl_w_ext                                           = int(0x87D8)
	gl_negative_x_ext                                  = int(0x87D9)
	gl_negative_y_ext                                  = int(0x87DA)
	gl_negative_z_ext                                  = int(0x87DB)
	gl_negative_w_ext                                  = int(0x87DC)
	gl_zero_ext                                        = int(0x87DD)
	gl_one_ext                                         = int(0x87DE)
	gl_negative_one_ext                                = int(0x87DF)
	gl_normalized_range_ext                            = int(0x87E0)
	gl_full_range_ext                                  = int(0x87E1)
	gl_current_vertex_ext                              = int(0x87E2)
	gl_mvp_matrix_ext                                  = int(0x87E3)
	gl_variant_value_ext                               = int(0x87E4)
	gl_variant_datatype_ext                            = int(0x87E5)
	gl_variant_array_stride_ext                        = int(0x87E6)
	gl_variant_array_type_ext                          = int(0x87E7)
	gl_variant_array_ext                               = int(0x87E8)
	gl_variant_array_pointer_ext                       = int(0x87E9)
	gl_invariant_value_ext                             = int(0x87EA)
	gl_invariant_datatype_ext                          = int(0x87EB)
	gl_local_constant_value_ext                        = int(0x87EC)
	gl_local_constant_datatype_ext                     = int(0x87ED)
	gl_atc_rgba_interpolated_alpha_amd                 = int(0x87EE)
	gl_pn_triangles_ati                                = int(0x87F0)
	gl_max_pn_triangles_tesselation_level_ati          = int(0x87F1)
	gl_pn_triangles_point_mode_ati                     = int(0x87F2)
	gl_pn_triangles_normal_mode_ati                    = int(0x87F3)
	gl_pn_triangles_tesselation_level_ati              = int(0x87F4)
	gl_pn_triangles_point_mode_linear_ati              = int(0x87F5)
	gl_pn_triangles_point_mode_cubic_ati               = int(0x87F6)
	gl_pn_triangles_normal_mode_linear_ati             = int(0x87F7)
	gl_pn_triangles_normal_mode_quadratic_ati          = int(0x87F8)
	gl_3dc_x_amd                                       = int(0x87F9)
	gl_3dc_xy_amd                                      = int(0x87FA)
	gl_vbo_free_memory_ati                             = int(0x87FB)
	gl_texture_free_memory_ati                         = int(0x87FC)
	gl_renderbuffer_free_memory_ati                    = int(0x87FD)
	gl_num_program_binary_formats                      = int(0x87FE)
	gl_num_program_binary_formats_oes                  = int(0x87FE)
	gl_program_binary_formats                          = int(0x87FF)
	gl_program_binary_formats_oes                      = int(0x87FF)
	gl_stencil_back_func                               = int(0x8800)
	gl_stencil_back_func_ati                           = int(0x8800)
	gl_stencil_back_fail                               = int(0x8801)
	gl_stencil_back_fail_ati                           = int(0x8801)
	gl_stencil_back_pass_depth_fail                    = int(0x8802)
	gl_stencil_back_pass_depth_fail_ati                = int(0x8802)
	gl_stencil_back_pass_depth_pass                    = int(0x8803)
	gl_stencil_back_pass_depth_pass_ati                = int(0x8803)
	gl_fragment_program_arb                            = int(0x8804)
	gl_program_alu_instructions_arb                    = int(0x8805)
	gl_program_tex_instructions_arb                    = int(0x8806)
	gl_program_tex_indirections_arb                    = int(0x8807)
	gl_program_native_alu_instructions_arb             = int(0x8808)
	gl_program_native_tex_instructions_arb             = int(0x8809)
	gl_program_native_tex_indirections_arb             = int(0x880A)
	gl_max_program_alu_instructions_arb                = int(0x880B)
	gl_max_program_tex_instructions_arb                = int(0x880C)
	gl_max_program_tex_indirections_arb                = int(0x880D)
	gl_max_program_native_alu_instructions_arb         = int(0x880E)
	gl_max_program_native_tex_instructions_arb         = int(0x880F)
	gl_max_program_native_tex_indirections_arb         = int(0x8810)
	gl_rgba32f                                         = int(0x8814)
	gl_rgba32f_arb                                     = int(0x8814)
	gl_rgba32f_ext                                     = int(0x8814)
	gl_rgba_float32_apple                              = int(0x8814)
	gl_rgba_float32_ati                                = int(0x8814)
	gl_rgb32f                                          = int(0x8815)
	gl_rgb32f_arb                                      = int(0x8815)
	gl_rgb32f_ext                                      = int(0x8815)
	gl_rgb_float32_apple                               = int(0x8815)
	gl_rgb_float32_ati                                 = int(0x8815)
	gl_alpha32f_arb                                    = int(0x8816)
	gl_alpha32f_ext                                    = int(0x8816)
	gl_alpha_float32_apple                             = int(0x8816)
	gl_alpha_float32_ati                               = int(0x8816)
	gl_intensity32f_arb                                = int(0x8817)
	gl_intensity_float32_apple                         = int(0x8817)
	gl_intensity_float32_ati                           = int(0x8817)
	gl_luminance32f_arb                                = int(0x8818)
	gl_luminance32f_ext                                = int(0x8818)
	gl_luminance_float32_apple                         = int(0x8818)
	gl_luminance_float32_ati                           = int(0x8818)
	gl_luminance_alpha32f_arb                          = int(0x8819)
	gl_luminance_alpha32f_ext                          = int(0x8819)
	gl_luminance_alpha_float32_apple                   = int(0x8819)
	gl_luminance_alpha_float32_ati                     = int(0x8819)
	gl_rgba16f                                         = int(0x881A)
	gl_rgba16f_arb                                     = int(0x881A)
	gl_rgba16f_ext                                     = int(0x881A)
	gl_rgba_float16_apple                              = int(0x881A)
	gl_rgba_float16_ati                                = int(0x881A)
	gl_rgb16f                                          = int(0x881B)
	gl_rgb16f_arb                                      = int(0x881B)
	gl_rgb16f_ext                                      = int(0x881B)
	gl_rgb_float16_apple                               = int(0x881B)
	gl_rgb_float16_ati                                 = int(0x881B)
	gl_alpha16f_arb                                    = int(0x881C)
	gl_alpha16f_ext                                    = int(0x881C)
	gl_alpha_float16_apple                             = int(0x881C)
	gl_alpha_float16_ati                               = int(0x881C)
	gl_intensity16f_arb                                = int(0x881D)
	gl_intensity_float16_apple                         = int(0x881D)
	gl_intensity_float16_ati                           = int(0x881D)
	gl_luminance16f_arb                                = int(0x881E)
	gl_luminance16f_ext                                = int(0x881E)
	gl_luminance_float16_apple                         = int(0x881E)
	gl_luminance_float16_ati                           = int(0x881E)
	gl_luminance_alpha16f_arb                          = int(0x881F)
	gl_luminance_alpha16f_ext                          = int(0x881F)
	gl_luminance_alpha_float16_apple                   = int(0x881F)
	gl_luminance_alpha_float16_ati                     = int(0x881F)
	gl_rgba_float_mode_arb                             = int(0x8820)
	gl_rgba_float_mode_ati                             = int(0x8820)
	gl_writeonly_rendering_qcom                        = int(0x8823)
	gl_max_draw_buffers                                = int(0x8824)
	gl_max_draw_buffers_arb                            = int(0x8824)
	gl_max_draw_buffers_ati                            = int(0x8824)
	gl_max_draw_buffers_ext                            = int(0x8824)
	gl_max_draw_buffers_nv                             = int(0x8824)
	gl_draw_buffer0                                    = int(0x8825)
	gl_draw_buffer0_arb                                = int(0x8825)
	gl_draw_buffer0_ati                                = int(0x8825)
	gl_draw_buffer0_ext                                = int(0x8825)
	gl_draw_buffer0_nv                                 = int(0x8825)
	gl_draw_buffer1                                    = int(0x8826)
	gl_draw_buffer1_arb                                = int(0x8826)
	gl_draw_buffer1_ati                                = int(0x8826)
	gl_draw_buffer1_ext                                = int(0x8826)
	gl_draw_buffer1_nv                                 = int(0x8826)
	gl_draw_buffer2                                    = int(0x8827)
	gl_draw_buffer2_arb                                = int(0x8827)
	gl_draw_buffer2_ati                                = int(0x8827)
	gl_draw_buffer2_ext                                = int(0x8827)
	gl_draw_buffer2_nv                                 = int(0x8827)
	gl_draw_buffer3                                    = int(0x8828)
	gl_draw_buffer3_arb                                = int(0x8828)
	gl_draw_buffer3_ati                                = int(0x8828)
	gl_draw_buffer3_ext                                = int(0x8828)
	gl_draw_buffer3_nv                                 = int(0x8828)
	gl_draw_buffer4                                    = int(0x8829)
	gl_draw_buffer4_arb                                = int(0x8829)
	gl_draw_buffer4_ati                                = int(0x8829)
	gl_draw_buffer4_ext                                = int(0x8829)
	gl_draw_buffer4_nv                                 = int(0x8829)
	gl_draw_buffer5                                    = int(0x882A)
	gl_draw_buffer5_arb                                = int(0x882A)
	gl_draw_buffer5_ati                                = int(0x882A)
	gl_draw_buffer5_ext                                = int(0x882A)
	gl_draw_buffer5_nv                                 = int(0x882A)
	gl_draw_buffer6                                    = int(0x882B)
	gl_draw_buffer6_arb                                = int(0x882B)
	gl_draw_buffer6_ati                                = int(0x882B)
	gl_draw_buffer6_ext                                = int(0x882B)
	gl_draw_buffer6_nv                                 = int(0x882B)
	gl_draw_buffer7                                    = int(0x882C)
	gl_draw_buffer7_arb                                = int(0x882C)
	gl_draw_buffer7_ati                                = int(0x882C)
	gl_draw_buffer7_ext                                = int(0x882C)
	gl_draw_buffer7_nv                                 = int(0x882C)
	gl_draw_buffer8                                    = int(0x882D)
	gl_draw_buffer8_arb                                = int(0x882D)
	gl_draw_buffer8_ati                                = int(0x882D)
	gl_draw_buffer8_ext                                = int(0x882D)
	gl_draw_buffer8_nv                                 = int(0x882D)
	gl_draw_buffer9                                    = int(0x882E)
	gl_draw_buffer9_arb                                = int(0x882E)
	gl_draw_buffer9_ati                                = int(0x882E)
	gl_draw_buffer9_ext                                = int(0x882E)
	gl_draw_buffer9_nv                                 = int(0x882E)
	gl_draw_buffer10                                   = int(0x882F)
	gl_draw_buffer10_arb                               = int(0x882F)
	gl_draw_buffer10_ati                               = int(0x882F)
	gl_draw_buffer10_ext                               = int(0x882F)
	gl_draw_buffer10_nv                                = int(0x882F)
	gl_draw_buffer11                                   = int(0x8830)
	gl_draw_buffer11_arb                               = int(0x8830)
	gl_draw_buffer11_ati                               = int(0x8830)
	gl_draw_buffer11_ext                               = int(0x8830)
	gl_draw_buffer11_nv                                = int(0x8830)
	gl_draw_buffer12                                   = int(0x8831)
	gl_draw_buffer12_arb                               = int(0x8831)
	gl_draw_buffer12_ati                               = int(0x8831)
	gl_draw_buffer12_ext                               = int(0x8831)
	gl_draw_buffer12_nv                                = int(0x8831)
	gl_draw_buffer13                                   = int(0x8832)
	gl_draw_buffer13_arb                               = int(0x8832)
	gl_draw_buffer13_ati                               = int(0x8832)
	gl_draw_buffer13_ext                               = int(0x8832)
	gl_draw_buffer13_nv                                = int(0x8832)
	gl_draw_buffer14                                   = int(0x8833)
	gl_draw_buffer14_arb                               = int(0x8833)
	gl_draw_buffer14_ati                               = int(0x8833)
	gl_draw_buffer14_ext                               = int(0x8833)
	gl_draw_buffer14_nv                                = int(0x8833)
	gl_draw_buffer15                                   = int(0x8834)
	gl_draw_buffer15_arb                               = int(0x8834)
	gl_draw_buffer15_ati                               = int(0x8834)
	gl_draw_buffer15_ext                               = int(0x8834)
	gl_draw_buffer15_nv                                = int(0x8834)
	gl_color_clear_unclamped_value_ati                 = int(0x8835)
	gl_compressed_luminance_alpha_3dc_ati              = int(0x8837)
	gl_blend_equation_alpha                            = int(0x883D)
	gl_blend_equation_alpha_ext                        = int(0x883D)
	gl_blend_equation_alpha_oes                        = int(0x883D)
	gl_subsample_distance_amd                          = int(0x883F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8840" end="0x884F" vendor="ARB" |>
pub const (
	gl_matrix_palette_arb                 = int(0x8840)
	gl_matrix_palette_oes                 = int(0x8840)
	gl_max_matrix_palette_stack_depth_arb = int(0x8841)
	gl_max_palette_matrices_arb           = int(0x8842)
	gl_max_palette_matrices_oes           = int(0x8842)
	gl_current_palette_matrix_arb         = int(0x8843)
	gl_current_palette_matrix_oes         = int(0x8843)
	gl_matrix_index_array_arb             = int(0x8844)
	gl_matrix_index_array_oes             = int(0x8844)
	gl_current_matrix_index_arb           = int(0x8845)
	gl_matrix_index_array_size_arb        = int(0x8846)
	gl_matrix_index_array_size_oes        = int(0x8846)
	gl_matrix_index_array_type_arb        = int(0x8847)
	gl_matrix_index_array_type_oes        = int(0x8847)
	gl_matrix_index_array_stride_arb      = int(0x8848)
	gl_matrix_index_array_stride_oes      = int(0x8848)
	gl_matrix_index_array_pointer_arb     = int(0x8849)
	gl_matrix_index_array_pointer_oes     = int(0x8849)
	gl_texture_depth_size                 = int(0x884A)
	gl_texture_depth_size_arb             = int(0x884A)
	gl_depth_texture_mode                 = int(0x884B)
	gl_depth_texture_mode_arb             = int(0x884B)
	gl_texture_compare_mode               = int(0x884C)
	gl_texture_compare_mode_arb           = int(0x884C)
	gl_texture_compare_mode_ext           = int(0x884C)
	gl_texture_compare_func               = int(0x884D)
	gl_texture_compare_func_arb           = int(0x884D)
	gl_texture_compare_func_ext           = int(0x884D)
	gl_compare_r_to_texture               = int(0x884E)
	gl_compare_r_to_texture_arb           = int(0x884E)
	gl_compare_ref_depth_to_texture_ext   = int(0x884E)
	gl_compare_ref_to_texture             = int(0x884E)
	gl_compare_ref_to_texture_ext         = int(0x884E)
	gl_texture_cube_map_seamless          = int(0x884F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8850" end="0x891F" vendor="NV" |>
pub const (
	gl_offset_projective_texture_2d_nv              = int(0x8850)
	gl_offset_projective_texture_2d_scale_nv        = int(0x8851)
	gl_offset_projective_texture_rectangle_nv       = int(0x8852)
	gl_offset_projective_texture_rectangle_scale_nv = int(0x8853)
	gl_offset_hilo_texture_2d_nv                    = int(0x8854)
	gl_offset_hilo_texture_rectangle_nv             = int(0x8855)
	gl_offset_hilo_projective_texture_2d_nv         = int(0x8856)
	gl_offset_hilo_projective_texture_rectangle_nv  = int(0x8857)
	gl_dependent_hilo_texture_2d_nv                 = int(0x8858)
	gl_dependent_rgb_texture_3d_nv                  = int(0x8859)
	gl_dependent_rgb_texture_cube_map_nv            = int(0x885A)
	gl_dot_product_pass_through_nv                  = int(0x885B)
	gl_dot_product_texture_1d_nv                    = int(0x885C)
	gl_dot_product_affine_depth_replace_nv          = int(0x885D)
	gl_hilo8_nv                                     = int(0x885E)
	gl_signed_hilo8_nv                              = int(0x885F)
	gl_force_blue_to_one_nv                         = int(0x8860)
	gl_point_sprite                                 = int(0x8861)
	gl_point_sprite_arb                             = int(0x8861)
	gl_point_sprite_nv                              = int(0x8861)
	gl_point_sprite_oes                             = int(0x8861)
	gl_coord_replace                                = int(0x8862)
	gl_coord_replace_arb                            = int(0x8862)
	gl_coord_replace_nv                             = int(0x8862)
	gl_coord_replace_oes                            = int(0x8862)
	gl_point_sprite_r_mode_nv                       = int(0x8863)
	gl_pixel_counter_bits_nv                        = int(0x8864)
	gl_query_counter_bits                           = int(0x8864)
	gl_query_counter_bits_arb                       = int(0x8864)
	gl_query_counter_bits_ext                       = int(0x8864)
	gl_current_occlusion_query_id_nv                = int(0x8865)
	gl_current_query                                = int(0x8865)
	gl_current_query_arb                            = int(0x8865)
	gl_current_query_ext                            = int(0x8865)
	gl_pixel_count_nv                               = int(0x8866)
	gl_query_result                                 = int(0x8866)
	gl_query_result_arb                             = int(0x8866)
	gl_query_result_ext                             = int(0x8866)
	gl_pixel_count_available_nv                     = int(0x8867)
	gl_query_result_available                       = int(0x8867)
	gl_query_result_available_arb                   = int(0x8867)
	gl_query_result_available_ext                   = int(0x8867)
	gl_max_fragment_program_local_parameters_nv     = int(0x8868)
	gl_max_vertex_attribs                           = int(0x8869)
	gl_max_vertex_attribs_arb                       = int(0x8869)
	gl_vertex_attrib_array_normalized               = int(0x886A)
	gl_vertex_attrib_array_normalized_arb           = int(0x886A)
	gl_max_tess_control_input_components            = int(0x886C)
	gl_max_tess_control_input_components_ext        = int(0x886C)
	gl_max_tess_control_input_components_oes        = int(0x886C)
	gl_max_tess_evaluation_input_components         = int(0x886D)
	gl_max_tess_evaluation_input_components_ext     = int(0x886D)
	gl_max_tess_evaluation_input_components_oes     = int(0x886D)
	gl_depth_stencil_to_rgba_nv                     = int(0x886E)
	gl_depth_stencil_to_bgra_nv                     = int(0x886F)
	gl_fragment_program_nv                          = int(0x8870)
	gl_max_texture_coords                           = int(0x8871)
	gl_max_texture_coords_arb                       = int(0x8871)
	gl_max_texture_coords_nv                        = int(0x8871)
	gl_max_texture_image_units                      = int(0x8872)
	gl_max_texture_image_units_arb                  = int(0x8872)
	gl_max_texture_image_units_nv                   = int(0x8872)
	gl_fragment_program_binding_nv                  = int(0x8873)
	gl_program_error_string_arb                     = int(0x8874)
	gl_program_error_string_nv                      = int(0x8874)
	gl_program_format_ascii_arb                     = int(0x8875)
	gl_program_format_arb                           = int(0x8876)
	gl_write_pixel_data_range_nv                    = int(0x8878)
	gl_read_pixel_data_range_nv                     = int(0x8879)
	gl_write_pixel_data_range_length_nv             = int(0x887A)
	gl_read_pixel_data_range_length_nv              = int(0x887B)
	gl_write_pixel_data_range_pointer_nv            = int(0x887C)
	gl_read_pixel_data_range_pointer_nv             = int(0x887D)
	gl_geometry_shader_invocations                  = int(0x887F)
	gl_geometry_shader_invocations_ext              = int(0x887F)
	gl_geometry_shader_invocations_oes              = int(0x887F)
	gl_float_r_nv                                   = int(0x8880)
	gl_float_rg_nv                                  = int(0x8881)
	gl_float_rgb_nv                                 = int(0x8882)
	gl_float_rgba_nv                                = int(0x8883)
	gl_float_r16_nv                                 = int(0x8884)
	gl_float_r32_nv                                 = int(0x8885)
	gl_float_rg16_nv                                = int(0x8886)
	gl_float_rg32_nv                                = int(0x8887)
	gl_float_rgb16_nv                               = int(0x8888)
	gl_float_rgb32_nv                               = int(0x8889)
	gl_float_rgba16_nv                              = int(0x888A)
	gl_float_rgba32_nv                              = int(0x888B)
	gl_texture_float_components_nv                  = int(0x888C)
	gl_float_clear_color_value_nv                   = int(0x888D)
	gl_float_rgba_mode_nv                           = int(0x888E)
	gl_texture_unsigned_remap_mode_nv               = int(0x888F)
	gl_depth_bounds_test_ext                        = int(0x8890)
	gl_depth_bounds_ext                             = int(0x8891)
	gl_array_buffer                                 = int(0x8892)
	gl_array_buffer_arb                             = int(0x8892)
	gl_element_array_buffer                         = int(0x8893)
	gl_element_array_buffer_arb                     = int(0x8893)
	gl_array_buffer_binding                         = int(0x8894)
	gl_array_buffer_binding_arb                     = int(0x8894)
	gl_element_array_buffer_binding                 = int(0x8895)
	gl_element_array_buffer_binding_arb             = int(0x8895)
	gl_vertex_array_buffer_binding                  = int(0x8896)
	gl_vertex_array_buffer_binding_arb              = int(0x8896)
	gl_normal_array_buffer_binding                  = int(0x8897)
	gl_normal_array_buffer_binding_arb              = int(0x8897)
	gl_color_array_buffer_binding                   = int(0x8898)
	gl_color_array_buffer_binding_arb               = int(0x8898)
	gl_index_array_buffer_binding                   = int(0x8899)
	gl_index_array_buffer_binding_arb               = int(0x8899)
	gl_texture_coord_array_buffer_binding           = int(0x889A)
	gl_texture_coord_array_buffer_binding_arb       = int(0x889A)
	gl_edge_flag_array_buffer_binding               = int(0x889B)
	gl_edge_flag_array_buffer_binding_arb           = int(0x889B)
	gl_secondary_color_array_buffer_binding         = int(0x889C)
	gl_secondary_color_array_buffer_binding_arb     = int(0x889C)
	gl_fog_coordinate_array_buffer_binding_arb      = int(0x889D)
	gl_fog_coordinate_array_buffer_binding          = int(0x889D)
	gl_fog_coord_array_buffer_binding               = int(0x889D)
	gl_weight_array_buffer_binding                  = int(0x889E)
	gl_weight_array_buffer_binding_arb              = int(0x889E)
	gl_weight_array_buffer_binding_oes              = int(0x889E)
	gl_vertex_attrib_array_buffer_binding           = int(0x889F)
	gl_vertex_attrib_array_buffer_binding_arb       = int(0x889F)
	gl_program_instructions_arb                     = int(0x88A0)
	gl_max_program_instructions_arb                 = int(0x88A1)
	gl_program_native_instructions_arb              = int(0x88A2)
	gl_max_program_native_instructions_arb          = int(0x88A3)
	gl_program_temporaries_arb                      = int(0x88A4)
	gl_max_program_temporaries_arb                  = int(0x88A5)
	gl_program_native_temporaries_arb               = int(0x88A6)
	gl_max_program_native_temporaries_arb           = int(0x88A7)
	gl_program_parameters_arb                       = int(0x88A8)
	gl_max_program_parameters_arb                   = int(0x88A9)
	gl_program_native_parameters_arb                = int(0x88AA)
	gl_max_program_native_parameters_arb            = int(0x88AB)
	gl_program_attribs_arb                          = int(0x88AC)
	gl_max_program_attribs_arb                      = int(0x88AD)
	gl_program_native_attribs_arb                   = int(0x88AE)
	gl_max_program_native_attribs_arb               = int(0x88AF)
	gl_program_address_registers_arb                = int(0x88B0)
	gl_max_program_address_registers_arb            = int(0x88B1)
	gl_program_native_address_registers_arb         = int(0x88B2)
	gl_max_program_native_address_registers_arb     = int(0x88B3)
	gl_max_program_local_parameters_arb             = int(0x88B4)
	gl_max_program_env_parameters_arb               = int(0x88B5)
	gl_program_under_native_limits_arb              = int(0x88B6)
	gl_transpose_current_matrix_arb                 = int(0x88B7)
	gl_read_only                                    = int(0x88B8)
	gl_read_only_arb                                = int(0x88B8)
	gl_write_only                                   = int(0x88B9)
	gl_write_only_arb                               = int(0x88B9)
	gl_write_only_oes                               = int(0x88B9)
	gl_read_write                                   = int(0x88BA)
	gl_read_write_arb                               = int(0x88BA)
	gl_buffer_access                                = int(0x88BB)
	gl_buffer_access_arb                            = int(0x88BB)
	gl_buffer_access_oes                            = int(0x88BB)
	gl_buffer_mapped                                = int(0x88BC)
	gl_buffer_mapped_arb                            = int(0x88BC)
	gl_buffer_mapped_oes                            = int(0x88BC)
	gl_buffer_map_pointer                           = int(0x88BD)
	gl_buffer_map_pointer_arb                       = int(0x88BD)
	gl_buffer_map_pointer_oes                       = int(0x88BD)
	gl_write_discard_nv                             = int(0x88BE)
	gl_time_elapsed                                 = int(0x88BF)
	gl_time_elapsed_ext                             = int(0x88BF)
	gl_matrix0_arb                                  = int(0x88C0)
	gl_matrix1_arb                                  = int(0x88C1)
	gl_matrix2_arb                                  = int(0x88C2)
	gl_matrix3_arb                                  = int(0x88C3)
	gl_matrix4_arb                                  = int(0x88C4)
	gl_matrix5_arb                                  = int(0x88C5)
	gl_matrix6_arb                                  = int(0x88C6)
	gl_matrix7_arb                                  = int(0x88C7)
	gl_matrix8_arb                                  = int(0x88C8)
	gl_matrix9_arb                                  = int(0x88C9)
	gl_matrix10_arb                                 = int(0x88CA)
	gl_matrix11_arb                                 = int(0x88CB)
	gl_matrix12_arb                                 = int(0x88CC)
	gl_matrix13_arb                                 = int(0x88CD)
	gl_matrix14_arb                                 = int(0x88CE)
	gl_matrix15_arb                                 = int(0x88CF)
	gl_matrix16_arb                                 = int(0x88D0)
	gl_matrix17_arb                                 = int(0x88D1)
	gl_matrix18_arb                                 = int(0x88D2)
	gl_matrix19_arb                                 = int(0x88D3)
	gl_matrix20_arb                                 = int(0x88D4)
	gl_matrix21_arb                                 = int(0x88D5)
	gl_matrix22_arb                                 = int(0x88D6)
	gl_matrix23_arb                                 = int(0x88D7)
	gl_matrix24_arb                                 = int(0x88D8)
	gl_matrix25_arb                                 = int(0x88D9)
	gl_matrix26_arb                                 = int(0x88DA)
	gl_matrix27_arb                                 = int(0x88DB)
	gl_matrix28_arb                                 = int(0x88DC)
	gl_matrix29_arb                                 = int(0x88DD)
	gl_matrix30_arb                                 = int(0x88DE)
	gl_matrix31_arb                                 = int(0x88DF)
	gl_stream_draw                                  = int(0x88E0)
	gl_stream_draw_arb                              = int(0x88E0)
	gl_stream_read                                  = int(0x88E1)
	gl_stream_read_arb                              = int(0x88E1)
	gl_stream_copy                                  = int(0x88E2)
	gl_stream_copy_arb                              = int(0x88E2)
	gl_static_draw                                  = int(0x88E4)
	gl_static_draw_arb                              = int(0x88E4)
	gl_static_read                                  = int(0x88E5)
	gl_static_read_arb                              = int(0x88E5)
	gl_static_copy                                  = int(0x88E6)
	gl_static_copy_arb                              = int(0x88E6)
	gl_dynamic_draw                                 = int(0x88E8)
	gl_dynamic_draw_arb                             = int(0x88E8)
	gl_dynamic_read                                 = int(0x88E9)
	gl_dynamic_read_arb                             = int(0x88E9)
	gl_dynamic_copy                                 = int(0x88EA)
	gl_dynamic_copy_arb                             = int(0x88EA)
	gl_pixel_pack_buffer                            = int(0x88EB)
	gl_pixel_pack_buffer_arb                        = int(0x88EB)
	gl_pixel_pack_buffer_ext                        = int(0x88EB)
	gl_pixel_pack_buffer_nv                         = int(0x88EB)
	gl_pixel_unpack_buffer                          = int(0x88EC)
	gl_pixel_unpack_buffer_arb                      = int(0x88EC)
	gl_pixel_unpack_buffer_ext                      = int(0x88EC)
	gl_pixel_unpack_buffer_nv                       = int(0x88EC)
	gl_pixel_pack_buffer_binding                    = int(0x88ED)
	gl_pixel_pack_buffer_binding_arb                = int(0x88ED)
	gl_pixel_pack_buffer_binding_ext                = int(0x88ED)
	gl_pixel_pack_buffer_binding_nv                 = int(0x88ED)
	gl_etc1_srgb8_nv                                = int(0x88EE)
	gl_pixel_unpack_buffer_binding                  = int(0x88EF)
	gl_pixel_unpack_buffer_binding_arb              = int(0x88EF)
	gl_pixel_unpack_buffer_binding_ext              = int(0x88EF)
	gl_pixel_unpack_buffer_binding_nv               = int(0x88EF)
	gl_depth24_stencil8                             = int(0x88F0)
	gl_depth24_stencil8_ext                         = int(0x88F0)
	gl_depth24_stencil8_oes                         = int(0x88F0)
	gl_texture_stencil_size                         = int(0x88F1)
	gl_texture_stencil_size_ext                     = int(0x88F1)
	gl_stencil_tag_bits_ext                         = int(0x88F2)
	gl_stencil_clear_tag_value_ext                  = int(0x88F3)
	gl_max_program_exec_instructions_nv             = int(0x88F4)
	gl_max_program_call_depth_nv                    = int(0x88F5)
	gl_max_program_if_depth_nv                      = int(0x88F6)
	gl_max_program_loop_depth_nv                    = int(0x88F7)
	gl_max_program_loop_count_nv                    = int(0x88F8)
	gl_src1_color                                   = int(0x88F9)
	gl_src1_color_ext                               = int(0x88F9)
	gl_one_minus_src1_color                         = int(0x88FA)
	gl_one_minus_src1_color_ext                     = int(0x88FA)
	gl_one_minus_src1_alpha                         = int(0x88FB)
	gl_one_minus_src1_alpha_ext                     = int(0x88FB)
	gl_max_dual_source_draw_buffers                 = int(0x88FC)
	gl_max_dual_source_draw_buffers_ext             = int(0x88FC)
	gl_vertex_attrib_array_integer                  = int(0x88FD)
	gl_vertex_attrib_array_integer_ext              = int(0x88FD)
	gl_vertex_attrib_array_integer_nv               = int(0x88FD)
	gl_vertex_attrib_array_divisor                  = int(0x88FE)
	gl_vertex_attrib_array_divisor_angle            = int(0x88FE)
	gl_vertex_attrib_array_divisor_arb              = int(0x88FE)
	gl_vertex_attrib_array_divisor_ext              = int(0x88FE)
	gl_vertex_attrib_array_divisor_nv               = int(0x88FE)
	gl_max_array_texture_layers                     = int(0x88FF)
	gl_max_array_texture_layers_ext                 = int(0x88FF)
	gl_min_program_texel_offset                     = int(0x8904)
	gl_min_program_texel_offset_ext                 = int(0x8904)
	gl_min_program_texel_offset_nv                  = int(0x8904)
	gl_max_program_texel_offset                     = int(0x8905)
	gl_max_program_texel_offset_ext                 = int(0x8905)
	gl_max_program_texel_offset_nv                  = int(0x8905)
	gl_program_attrib_components_nv                 = int(0x8906)
	gl_program_result_components_nv                 = int(0x8907)
	gl_max_program_attrib_components_nv             = int(0x8908)
	gl_max_program_result_components_nv             = int(0x8909)
	gl_stencil_test_two_side_ext                    = int(0x8910)
	gl_active_stencil_face_ext                      = int(0x8911)
	gl_mirror_clamp_to_border_ext                   = int(0x8912)
	gl_samples_passed                               = int(0x8914)
	gl_samples_passed_arb                           = int(0x8914)
	gl_geometry_vertices_out                        = int(0x8916)
	gl_geometry_linked_vertices_out_ext             = int(0x8916)
	gl_geometry_linked_vertices_out_oes             = int(0x8916)
	gl_geometry_input_type                          = int(0x8917)
	gl_geometry_linked_input_type_ext               = int(0x8917)
	gl_geometry_linked_input_type_oes               = int(0x8917)
	gl_geometry_output_type                         = int(0x8918)
	gl_geometry_linked_output_type_ext              = int(0x8918)
	gl_geometry_linked_output_type_oes              = int(0x8918)
	gl_sampler_binding                              = int(0x8919)
	gl_clamp_vertex_color                           = int(0x891A)
	gl_clamp_vertex_color_arb                       = int(0x891A)
	gl_clamp_fragment_color                         = int(0x891B)
	gl_clamp_fragment_color_arb                     = int(0x891B)
	gl_clamp_read_color                             = int(0x891C)
	gl_clamp_read_color_arb                         = int(0x891C)
	gl_fixed_only                                   = int(0x891D)
	gl_fixed_only_arb                               = int(0x891D)
	gl_tess_control_program_nv                      = int(0x891E)
	gl_tess_evaluation_program_nv                   = int(0x891F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8920" end="0x897F" vendor="AMD" |>
pub const (
	gl_fragment_shader_ati                   = int(0x8920)
	gl_reg_0_ati                             = int(0x8921)
	gl_reg_1_ati                             = int(0x8922)
	gl_reg_2_ati                             = int(0x8923)
	gl_reg_3_ati                             = int(0x8924)
	gl_reg_4_ati                             = int(0x8925)
	gl_reg_5_ati                             = int(0x8926)
	gl_reg_6_ati                             = int(0x8927)
	gl_reg_7_ati                             = int(0x8928)
	gl_reg_8_ati                             = int(0x8929)
	gl_reg_9_ati                             = int(0x892A)
	gl_reg_10_ati                            = int(0x892B)
	gl_reg_11_ati                            = int(0x892C)
	gl_reg_12_ati                            = int(0x892D)
	gl_reg_13_ati                            = int(0x892E)
	gl_reg_14_ati                            = int(0x892F)
	gl_reg_15_ati                            = int(0x8930)
	gl_reg_16_ati                            = int(0x8931)
	gl_reg_17_ati                            = int(0x8932)
	gl_reg_18_ati                            = int(0x8933)
	gl_reg_19_ati                            = int(0x8934)
	gl_reg_20_ati                            = int(0x8935)
	gl_reg_21_ati                            = int(0x8936)
	gl_reg_22_ati                            = int(0x8937)
	gl_reg_23_ati                            = int(0x8938)
	gl_reg_24_ati                            = int(0x8939)
	gl_reg_25_ati                            = int(0x893A)
	gl_reg_26_ati                            = int(0x893B)
	gl_reg_27_ati                            = int(0x893C)
	gl_reg_28_ati                            = int(0x893D)
	gl_reg_29_ati                            = int(0x893E)
	gl_reg_30_ati                            = int(0x893F)
	gl_reg_31_ati                            = int(0x8940)
	gl_con_0_ati                             = int(0x8941)
	gl_con_1_ati                             = int(0x8942)
	gl_con_2_ati                             = int(0x8943)
	gl_con_3_ati                             = int(0x8944)
	gl_con_4_ati                             = int(0x8945)
	gl_con_5_ati                             = int(0x8946)
	gl_con_6_ati                             = int(0x8947)
	gl_con_7_ati                             = int(0x8948)
	gl_con_8_ati                             = int(0x8949)
	gl_con_9_ati                             = int(0x894A)
	gl_con_10_ati                            = int(0x894B)
	gl_con_11_ati                            = int(0x894C)
	gl_con_12_ati                            = int(0x894D)
	gl_con_13_ati                            = int(0x894E)
	gl_con_14_ati                            = int(0x894F)
	gl_con_15_ati                            = int(0x8950)
	gl_con_16_ati                            = int(0x8951)
	gl_con_17_ati                            = int(0x8952)
	gl_con_18_ati                            = int(0x8953)
	gl_con_19_ati                            = int(0x8954)
	gl_con_20_ati                            = int(0x8955)
	gl_con_21_ati                            = int(0x8956)
	gl_con_22_ati                            = int(0x8957)
	gl_con_23_ati                            = int(0x8958)
	gl_con_24_ati                            = int(0x8959)
	gl_con_25_ati                            = int(0x895A)
	gl_con_26_ati                            = int(0x895B)
	gl_con_27_ati                            = int(0x895C)
	gl_con_28_ati                            = int(0x895D)
	gl_con_29_ati                            = int(0x895E)
	gl_con_30_ati                            = int(0x895F)
	gl_con_31_ati                            = int(0x8960)
	gl_mov_ati                               = int(0x8961)
	gl_add_ati                               = int(0x8963)
	gl_mul_ati                               = int(0x8964)
	gl_sub_ati                               = int(0x8965)
	gl_dot3_ati                              = int(0x8966)
	gl_dot4_ati                              = int(0x8967)
	gl_mad_ati                               = int(0x8968)
	gl_lerp_ati                              = int(0x8969)
	gl_cnd_ati                               = int(0x896A)
	gl_cnd0_ati                              = int(0x896B)
	gl_dot2_add_ati                          = int(0x896C)
	gl_secondary_interpolator_ati            = int(0x896D)
	gl_num_fragment_registers_ati            = int(0x896E)
	gl_num_fragment_constants_ati            = int(0x896F)
	gl_num_passes_ati                        = int(0x8970)
	gl_num_instructions_per_pass_ati         = int(0x8971)
	gl_num_instructions_total_ati            = int(0x8972)
	gl_num_input_interpolator_components_ati = int(0x8973)
	gl_num_loopback_components_ati           = int(0x8974)
	gl_color_alpha_pairing_ati               = int(0x8975)
	gl_swizzle_str_ati                       = int(0x8976)
	gl_swizzle_stq_ati                       = int(0x8977)
	gl_swizzle_str_dr_ati                    = int(0x8978)
	gl_swizzle_stq_dq_ati                    = int(0x8979)
	gl_swizzle_strq_ati                      = int(0x897A)
	gl_swizzle_strq_dq_ati                   = int(0x897B)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8980" end="0x898F" vendor="OML" |>
pub const (
	gl_interlace_oml                           = int(0x8980)
	gl_interlace_read_oml                      = int(0x8981)
	gl_format_subsample_24_24_oml              = int(0x8982)
	gl_format_subsample_244_244_oml            = int(0x8983)
	gl_pack_resample_oml                       = int(0x8984)
	gl_unpack_resample_oml                     = int(0x8985)
	gl_resample_replicate_oml                  = int(0x8986)
	gl_resample_zero_fill_oml                  = int(0x8987)
	gl_resample_average_oml                    = int(0x8988)
	gl_resample_decimate_oml                   = int(0x8989)
	gl_point_size_array_type_oes               = int(0x898A)
	gl_point_size_array_stride_oes             = int(0x898B)
	gl_point_size_array_pointer_oes            = int(0x898C)
	gl_modelview_matrix_float_as_int_bits_oes  = int(0x898D)
	gl_projection_matrix_float_as_int_bits_oes = int(0x898E)
	gl_texture_matrix_float_as_int_bits_oes    = int(0x898F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8A00" end="0x8A7F" vendor="APPLE" |>
pub const (
	gl_vertex_attrib_map1_apple                     = int(0x8A00)
	gl_vertex_attrib_map2_apple                     = int(0x8A01)
	gl_vertex_attrib_map1_size_apple                = int(0x8A02)
	gl_vertex_attrib_map1_coeff_apple               = int(0x8A03)
	gl_vertex_attrib_map1_order_apple               = int(0x8A04)
	gl_vertex_attrib_map1_domain_apple              = int(0x8A05)
	gl_vertex_attrib_map2_size_apple                = int(0x8A06)
	gl_vertex_attrib_map2_coeff_apple               = int(0x8A07)
	gl_vertex_attrib_map2_order_apple               = int(0x8A08)
	gl_vertex_attrib_map2_domain_apple              = int(0x8A09)
	gl_draw_pixels_apple                            = int(0x8A0A)
	gl_fence_apple                                  = int(0x8A0B)
	gl_element_array_apple                          = int(0x8A0C)
	gl_element_array_type_apple                     = int(0x8A0D)
	gl_element_array_pointer_apple                  = int(0x8A0E)
	gl_color_float_apple                            = int(0x8A0F)
	gl_uniform_buffer                               = int(0x8A11)
	gl_buffer_serialized_modify_apple               = int(0x8A12)
	gl_buffer_flushing_unmap_apple                  = int(0x8A13)
	gl_aux_depth_stencil_apple                      = int(0x8A14)
	gl_pack_row_bytes_apple                         = int(0x8A15)
	gl_unpack_row_bytes_apple                       = int(0x8A16)
	gl_released_apple                               = int(0x8A19)
	gl_volatile_apple                               = int(0x8A1A)
	gl_retained_apple                               = int(0x8A1B)
	gl_undefined_apple                              = int(0x8A1C)
	gl_purgeable_apple                              = int(0x8A1D)
	gl_rgb_422_apple                                = int(0x8A1F)
	gl_uniform_buffer_binding                       = int(0x8A28)
	gl_uniform_buffer_start                         = int(0x8A29)
	gl_uniform_buffer_size                          = int(0x8A2A)
	gl_max_vertex_uniform_blocks                    = int(0x8A2B)
	gl_max_geometry_uniform_blocks                  = int(0x8A2C)
	gl_max_geometry_uniform_blocks_ext              = int(0x8A2C)
	gl_max_geometry_uniform_blocks_oes              = int(0x8A2C)
	gl_max_fragment_uniform_blocks                  = int(0x8A2D)
	gl_max_combined_uniform_blocks                  = int(0x8A2E)
	gl_max_uniform_buffer_bindings                  = int(0x8A2F)
	gl_max_uniform_block_size                       = int(0x8A30)
	gl_max_combined_vertex_uniform_components       = int(0x8A31)
	gl_max_combined_geometry_uniform_components     = int(0x8A32)
	gl_max_combined_geometry_uniform_components_ext = int(0x8A32)
	gl_max_combined_geometry_uniform_components_oes = int(0x8A32)
	gl_max_combined_fragment_uniform_components     = int(0x8A33)
	gl_uniform_buffer_offset_alignment              = int(0x8A34)
	gl_active_uniform_block_max_name_length         = int(0x8A35)
	gl_active_uniform_blocks                        = int(0x8A36)
	gl_uniform_type                                 = int(0x8A37)
	gl_uniform_size                                 = int(0x8A38)
	gl_uniform_name_length                          = int(0x8A39)
	gl_uniform_block_index                          = int(0x8A3A)
	gl_uniform_offset                               = int(0x8A3B)
	gl_uniform_array_stride                         = int(0x8A3C)
	gl_uniform_matrix_stride                        = int(0x8A3D)
	gl_uniform_is_row_major                         = int(0x8A3E)
	gl_uniform_block_binding                        = int(0x8A3F)
	gl_uniform_block_data_size                      = int(0x8A40)
	gl_uniform_block_name_length                    = int(0x8A41)
	gl_uniform_block_active_uniforms                = int(0x8A42)
	gl_uniform_block_active_uniform_indices         = int(0x8A43)
	gl_uniform_block_referenced_by_vertex_shader    = int(0x8A44)
	gl_uniform_block_referenced_by_geometry_shader  = int(0x8A45)
	gl_uniform_block_referenced_by_fragment_shader  = int(0x8A46)
	gl_texture_srgb_decode_ext                      = int(0x8A48)
	gl_decode_ext                                   = int(0x8A49)
	gl_skip_decode_ext                              = int(0x8A4A)
	gl_program_pipeline_object_ext                  = int(0x8A4F)
	gl_rgb_raw_422_apple                            = int(0x8A51)
	gl_fragment_shader_discards_samples_ext         = int(0x8A52)
	gl_sync_object_apple                            = int(0x8A53)
	gl_compressed_srgb_pvrtc_2bppv1_ext             = int(0x8A54)
	gl_compressed_srgb_pvrtc_4bppv1_ext             = int(0x8A55)
	gl_compressed_srgb_alpha_pvrtc_2bppv1_ext       = int(0x8A56)
	gl_compressed_srgb_alpha_pvrtc_4bppv1_ext       = int(0x8A57)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8B30" end="0x8B3F" group="ShaderType" vendor="ARB" |>
pub const (
	gl_fragment_shader     = int(0x8B30)
	gl_fragment_shader_arb = int(0x8B30)
	gl_vertex_shader       = int(0x8B31)
	gl_vertex_shader_arb   = int(0x8B31)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8B40" end="0x8B47" group="ContainerType" vendor="ARB" |>
pub const (
	gl_program_object_arb = int(0x8B40)
	gl_program_object_ext = int(0x8B40)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8B48" end="0x8B4F" vendor="ARB" |>
pub const (
	gl_shader_object_arb                    = int(0x8B48)
	gl_shader_object_ext                    = int(0x8B48)
	gl_max_fragment_uniform_components      = int(0x8B49)
	gl_max_fragment_uniform_components_arb  = int(0x8B49)
	gl_max_vertex_uniform_components        = int(0x8B4A)
	gl_max_vertex_uniform_components_arb    = int(0x8B4A)
	gl_max_varying_floats                   = int(0x8B4B)
	gl_max_varying_components               = int(0x8B4B)
	gl_max_varying_components_ext           = int(0x8B4B)
	gl_max_varying_floats_arb               = int(0x8B4B)
	gl_max_vertex_texture_image_units       = int(0x8B4C)
	gl_max_vertex_texture_image_units_arb   = int(0x8B4C)
	gl_max_combined_texture_image_units     = int(0x8B4D)
	gl_max_combined_texture_image_units_arb = int(0x8B4D)
	gl_object_type_arb                      = int(0x8B4E)
	gl_shader_type                          = int(0x8B4F)
	gl_object_subtype_arb                   = int(0x8B4F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8B50" end="0x8B7F" group="AttributeType" vendor="ARB" |>
pub const (
	gl_float_vec2                 = int(0x8B50)
	gl_float_vec2_arb             = int(0x8B50)
	gl_float_vec3                 = int(0x8B51)
	gl_float_vec3_arb             = int(0x8B51)
	gl_float_vec4                 = int(0x8B52)
	gl_float_vec4_arb             = int(0x8B52)
	gl_int_vec2                   = int(0x8B53)
	gl_int_vec2_arb               = int(0x8B53)
	gl_int_vec3                   = int(0x8B54)
	gl_int_vec3_arb               = int(0x8B54)
	gl_int_vec4                   = int(0x8B55)
	gl_int_vec4_arb               = int(0x8B55)
	gl_bool                       = int(0x8B56)
	gl_bool_arb                   = int(0x8B56)
	gl_bool_vec2                  = int(0x8B57)
	gl_bool_vec2_arb              = int(0x8B57)
	gl_bool_vec3                  = int(0x8B58)
	gl_bool_vec3_arb              = int(0x8B58)
	gl_bool_vec4                  = int(0x8B59)
	gl_bool_vec4_arb              = int(0x8B59)
	gl_float_mat2                 = int(0x8B5A)
	gl_float_mat2_arb             = int(0x8B5A)
	gl_float_mat3                 = int(0x8B5B)
	gl_float_mat3_arb             = int(0x8B5B)
	gl_float_mat4                 = int(0x8B5C)
	gl_float_mat4_arb             = int(0x8B5C)
	gl_sampler_1d                 = int(0x8B5D)
	gl_sampler_1d_arb             = int(0x8B5D)
	gl_sampler_2d                 = int(0x8B5E)
	gl_sampler_2d_arb             = int(0x8B5E)
	gl_sampler_3d                 = int(0x8B5F)
	gl_sampler_3d_arb             = int(0x8B5F)
	gl_sampler_3d_oes             = int(0x8B5F)
	gl_sampler_cube               = int(0x8B60)
	gl_sampler_cube_arb           = int(0x8B60)
	gl_sampler_1d_shadow          = int(0x8B61)
	gl_sampler_1d_shadow_arb      = int(0x8B61)
	gl_sampler_2d_shadow          = int(0x8B62)
	gl_sampler_2d_shadow_arb      = int(0x8B62)
	gl_sampler_2d_shadow_ext      = int(0x8B62)
	gl_sampler_2d_rect            = int(0x8B63)
	gl_sampler_2d_rect_arb        = int(0x8B63)
	gl_sampler_2d_rect_shadow     = int(0x8B64)
	gl_sampler_2d_rect_shadow_arb = int(0x8B64)
	gl_float_mat2x3               = int(0x8B65)
	gl_float_mat2x3_nv            = int(0x8B65)
	gl_float_mat2x4               = int(0x8B66)
	gl_float_mat2x4_nv            = int(0x8B66)
	gl_float_mat3x2               = int(0x8B67)
	gl_float_mat3x2_nv            = int(0x8B67)
	gl_float_mat3x4               = int(0x8B68)
	gl_float_mat3x4_nv            = int(0x8B68)
	gl_float_mat4x2               = int(0x8B69)
	gl_float_mat4x2_nv            = int(0x8B69)
	gl_float_mat4x3               = int(0x8B6A)
	gl_float_mat4x3_nv            = int(0x8B6A)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8B80" end="0x8B8F" vendor="ARB" |>
pub const (
	gl_delete_status                          = int(0x8B80)
	gl_object_delete_status_arb               = int(0x8B80)
	gl_compile_status                         = int(0x8B81)
	gl_object_compile_status_arb              = int(0x8B81)
	gl_link_status                            = int(0x8B82)
	gl_object_link_status_arb                 = int(0x8B82)
	gl_validate_status                        = int(0x8B83)
	gl_object_validate_status_arb             = int(0x8B83)
	gl_info_log_length                        = int(0x8B84)
	gl_object_info_log_length_arb             = int(0x8B84)
	gl_attached_shaders                       = int(0x8B85)
	gl_object_attached_objects_arb            = int(0x8B85)
	gl_active_uniforms                        = int(0x8B86)
	gl_object_active_uniforms_arb             = int(0x8B86)
	gl_active_uniform_max_length              = int(0x8B87)
	gl_object_active_uniform_max_length_arb   = int(0x8B87)
	gl_shader_source_length                   = int(0x8B88)
	gl_object_shader_source_length_arb        = int(0x8B88)
	gl_active_attributes                      = int(0x8B89)
	gl_object_active_attributes_arb           = int(0x8B89)
	gl_active_attribute_max_length            = int(0x8B8A)
	gl_object_active_attribute_max_length_arb = int(0x8B8A)
	gl_fragment_shader_derivative_hint        = int(0x8B8B)
	gl_fragment_shader_derivative_hint_arb    = int(0x8B8B)
	gl_fragment_shader_derivative_hint_oes    = int(0x8B8B)
	gl_shading_language_version               = int(0x8B8C)
	gl_shading_language_version_arb           = int(0x8B8C)
	gl_current_program                        = int(0x8B8D)
		// todo duplicate : gl_active_program_ext = int(0x8B8D)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8B90" end="0x8B9F" vendor="OES" |>
pub const (
	gl_palette4_rgb8_oes                     = int(0x8B90)
	gl_palette4_rgba8_oes                    = int(0x8B91)
	gl_palette4_r5_g6_b5_oes                 = int(0x8B92)
	gl_palette4_rgba4_oes                    = int(0x8B93)
	gl_palette4_rgb5_a1_oes                  = int(0x8B94)
	gl_palette8_rgb8_oes                     = int(0x8B95)
	gl_palette8_rgba8_oes                    = int(0x8B96)
	gl_palette8_r5_g6_b5_oes                 = int(0x8B97)
	gl_palette8_rgba4_oes                    = int(0x8B98)
	gl_palette8_rgb5_a1_oes                  = int(0x8B99)
	gl_implementation_color_read_type        = int(0x8B9A)
	gl_implementation_color_read_type_oes    = int(0x8B9A)
	gl_implementation_color_read_format      = int(0x8B9B)
	gl_implementation_color_read_format_oes  = int(0x8B9B)
	gl_point_size_array_oes                  = int(0x8B9C)
	gl_texture_crop_rect_oes                 = int(0x8B9D)
	gl_matrix_index_array_buffer_binding_oes = int(0x8B9E)
	gl_point_size_array_buffer_binding_oes   = int(0x8B9F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8BB0" end="0x8BBF" vendor="MESA" |>
pub const (
	gl_fragment_program_position_mesa      = int(0x8BB0)
	gl_fragment_program_callback_mesa      = int(0x8BB1)
	gl_fragment_program_callback_func_mesa = int(0x8BB2)
	gl_fragment_program_callback_data_mesa = int(0x8BB3)
	gl_vertex_program_position_mesa        = int(0x8BB4)
	gl_vertex_program_callback_mesa        = int(0x8BB5)
	gl_vertex_program_callback_func_mesa   = int(0x8BB6)
	gl_vertex_program_callback_data_mesa   = int(0x8BB7)
	gl_tile_raster_order_fixed_mesa        = int(0x8BB8)
	gl_tile_raster_order_increasing_x_mesa = int(0x8BB9)
	gl_tile_raster_order_increasing_y_mesa = int(0x8BBA)
	gl_framebuffer_flip_y_mesa             = int(0x8BBB)
	gl_framebuffer_flip_x_mesa             = int(0x8BBC)
	gl_framebuffer_swap_xy_mesa            = int(0x8BBD)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8BC0" end="0x8BFF" vendor="QCOM" comment="Reassigned from AMD to QCOM" |>
pub const (
	gl_counter_type_amd                             = int(0x8BC0)
	gl_counter_range_amd                            = int(0x8BC1)
	gl_unsigned_int64_amd                           = int(0x8BC2)
	gl_percentage_amd                               = int(0x8BC3)
	gl_perfmon_result_available_amd                 = int(0x8BC4)
	gl_perfmon_result_size_amd                      = int(0x8BC5)
	gl_perfmon_result_amd                           = int(0x8BC6)
	gl_texture_width_qcom                           = int(0x8BD2)
	gl_texture_height_qcom                          = int(0x8BD3)
	gl_texture_depth_qcom                           = int(0x8BD4)
	gl_texture_internal_format_qcom                 = int(0x8BD5)
	gl_texture_format_qcom                          = int(0x8BD6)
	gl_texture_type_qcom                            = int(0x8BD7)
	gl_texture_image_valid_qcom                     = int(0x8BD8)
	gl_texture_num_levels_qcom                      = int(0x8BD9)
	gl_texture_target_qcom                          = int(0x8BDA)
	gl_texture_object_valid_qcom                    = int(0x8BDB)
	gl_state_restore                                = int(0x8BDC)
	gl_sampler_external_2d_y2y_ext                  = int(0x8BE7)
	gl_texture_protected_ext                        = int(0x8BFA)
	gl_texture_foveated_feature_bits_qcom           = int(0x8BFB)
	gl_texture_foveated_min_pixel_density_qcom      = int(0x8BFC)
	gl_texture_foveated_feature_query_qcom          = int(0x8BFD)
	gl_texture_foveated_num_focal_points_query_qcom = int(0x8BFE)
	gl_framebuffer_incomplete_foveation_qcom        = int(0x8BFF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8C00" end="0x8C0F" vendor="IMG" |>
pub const (
	gl_compressed_rgb_pvrtc_4bppv1_img  = int(0x8C00)
	gl_compressed_rgb_pvrtc_2bppv1_img  = int(0x8C01)
	gl_compressed_rgba_pvrtc_4bppv1_img = int(0x8C02)
	gl_compressed_rgba_pvrtc_2bppv1_img = int(0x8C03)
	gl_modulate_color_img               = int(0x8C04)
	gl_recip_add_signed_alpha_img       = int(0x8C05)
	gl_texture_alpha_modulate_img       = int(0x8C06)
	gl_factor_alpha_modulate_img        = int(0x8C07)
	gl_fragment_alpha_modulate_img      = int(0x8C08)
	gl_add_blend_img                    = int(0x8C09)
	gl_sgx_binary_img                   = int(0x8C0A)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8C10" end="0x8C8F" vendor="NV" comment="For Pat Brown" |>
pub const (
	gl_texture_red_type                                  = int(0x8C10)
	gl_texture_red_type_arb                              = int(0x8C10)
	gl_texture_green_type                                = int(0x8C11)
	gl_texture_green_type_arb                            = int(0x8C11)
	gl_texture_blue_type                                 = int(0x8C12)
	gl_texture_blue_type_arb                             = int(0x8C12)
	gl_texture_alpha_type                                = int(0x8C13)
	gl_texture_alpha_type_arb                            = int(0x8C13)
	gl_texture_luminance_type                            = int(0x8C14)
	gl_texture_luminance_type_arb                        = int(0x8C14)
	gl_texture_intensity_type                            = int(0x8C15)
	gl_texture_intensity_type_arb                        = int(0x8C15)
	gl_texture_depth_type                                = int(0x8C16)
	gl_texture_depth_type_arb                            = int(0x8C16)
	gl_unsigned_normalized                               = int(0x8C17)
	gl_unsigned_normalized_arb                           = int(0x8C17)
	gl_unsigned_normalized_ext                           = int(0x8C17)
	gl_texture_1d_array                                  = int(0x8C18)
	gl_texture_1d_array_ext                              = int(0x8C18)
	gl_proxy_texture_1d_array                            = int(0x8C19)
	gl_proxy_texture_1d_array_ext                        = int(0x8C19)
	gl_texture_2d_array                                  = int(0x8C1A)
	gl_texture_2d_array_ext                              = int(0x8C1A)
	gl_proxy_texture_2d_array                            = int(0x8C1B)
	gl_proxy_texture_2d_array_ext                        = int(0x8C1B)
	gl_texture_binding_1d_array                          = int(0x8C1C)
	gl_texture_binding_1d_array_ext                      = int(0x8C1C)
	gl_texture_binding_2d_array                          = int(0x8C1D)
	gl_texture_binding_2d_array_ext                      = int(0x8C1D)
	gl_geometry_program_nv                               = int(0x8C26)
	gl_max_program_output_vertices_nv                    = int(0x8C27)
	gl_max_program_total_output_components_nv            = int(0x8C28)
	gl_max_geometry_texture_image_units                  = int(0x8C29)
	gl_max_geometry_texture_image_units_arb              = int(0x8C29)
	gl_max_geometry_texture_image_units_ext              = int(0x8C29)
	gl_max_geometry_texture_image_units_oes              = int(0x8C29)
	gl_texture_buffer                                    = int(0x8C2A)
	gl_texture_buffer_arb                                = int(0x8C2A)
	gl_texture_buffer_ext                                = int(0x8C2A)
	gl_texture_buffer_oes                                = int(0x8C2A)
	gl_texture_buffer_binding                            = int(0x8C2A)
	gl_texture_buffer_binding_ext                        = int(0x8C2A)
	gl_texture_buffer_binding_oes                        = int(0x8C2A)
	gl_max_texture_buffer_size                           = int(0x8C2B)
	gl_max_texture_buffer_size_arb                       = int(0x8C2B)
	gl_max_texture_buffer_size_ext                       = int(0x8C2B)
	gl_max_texture_buffer_size_oes                       = int(0x8C2B)
	gl_texture_binding_buffer                            = int(0x8C2C)
	gl_texture_binding_buffer_arb                        = int(0x8C2C)
	gl_texture_binding_buffer_ext                        = int(0x8C2C)
	gl_texture_binding_buffer_oes                        = int(0x8C2C)
	gl_texture_buffer_data_store_binding                 = int(0x8C2D)
	gl_texture_buffer_data_store_binding_arb             = int(0x8C2D)
	gl_texture_buffer_data_store_binding_ext             = int(0x8C2D)
	gl_texture_buffer_data_store_binding_oes             = int(0x8C2D)
	gl_texture_buffer_format_arb                         = int(0x8C2E)
	gl_texture_buffer_format_ext                         = int(0x8C2E)
	gl_any_samples_passed                                = int(0x8C2F)
	gl_any_samples_passed_ext                            = int(0x8C2F)
	gl_sample_shading                                    = int(0x8C36)
	gl_sample_shading_arb                                = int(0x8C36)
	gl_sample_shading_oes                                = int(0x8C36)
	gl_min_sample_shading_value                          = int(0x8C37)
	gl_min_sample_shading_value_arb                      = int(0x8C37)
	gl_min_sample_shading_value_oes                      = int(0x8C37)
	gl_r11f_g11f_b10f                                    = int(0x8C3A)
	gl_r11f_g11f_b10f_apple                              = int(0x8C3A)
	gl_r11f_g11f_b10f_ext                                = int(0x8C3A)
	gl_unsigned_int_10f_11f_11f_rev                      = int(0x8C3B)
	gl_unsigned_int_10f_11f_11f_rev_apple                = int(0x8C3B)
	gl_unsigned_int_10f_11f_11f_rev_ext                  = int(0x8C3B)
	gl_rgba_signed_components_ext                        = int(0x8C3C)
	gl_rgb9_e5                                           = int(0x8C3D)
	gl_rgb9_e5_apple                                     = int(0x8C3D)
	gl_rgb9_e5_ext                                       = int(0x8C3D)
	gl_unsigned_int_5_9_9_9_rev                          = int(0x8C3E)
	gl_unsigned_int_5_9_9_9_rev_apple                    = int(0x8C3E)
	gl_unsigned_int_5_9_9_9_rev_ext                      = int(0x8C3E)
	gl_texture_shared_size                               = int(0x8C3F)
	gl_texture_shared_size_ext                           = int(0x8C3F)
	gl_srgb                                              = int(0x8C40)
	gl_srgb_ext                                          = int(0x8C40)
	gl_srgb8                                             = int(0x8C41)
	gl_srgb8_ext                                         = int(0x8C41)
	gl_srgb8_nv                                          = int(0x8C41)
	gl_srgb_alpha                                        = int(0x8C42)
	gl_srgb_alpha_ext                                    = int(0x8C42)
	gl_srgb8_alpha8                                      = int(0x8C43)
	gl_srgb8_alpha8_ext                                  = int(0x8C43)
	gl_sluminance_alpha                                  = int(0x8C44)
	gl_sluminance_alpha_ext                              = int(0x8C44)
	gl_sluminance_alpha_nv                               = int(0x8C44)
	gl_sluminance8_alpha8                                = int(0x8C45)
	gl_sluminance8_alpha8_ext                            = int(0x8C45)
	gl_sluminance8_alpha8_nv                             = int(0x8C45)
	gl_sluminance                                        = int(0x8C46)
	gl_sluminance_ext                                    = int(0x8C46)
	gl_sluminance_nv                                     = int(0x8C46)
	gl_sluminance8                                       = int(0x8C47)
	gl_sluminance8_ext                                   = int(0x8C47)
	gl_sluminance8_nv                                    = int(0x8C47)
	gl_compressed_srgb                                   = int(0x8C48)
	gl_compressed_srgb_ext                               = int(0x8C48)
	gl_compressed_srgb_alpha                             = int(0x8C49)
	gl_compressed_srgb_alpha_ext                         = int(0x8C49)
	gl_compressed_sluminance                             = int(0x8C4A)
	gl_compressed_sluminance_ext                         = int(0x8C4A)
	gl_compressed_sluminance_alpha                       = int(0x8C4B)
	gl_compressed_sluminance_alpha_ext                   = int(0x8C4B)
	gl_compressed_srgb_s3tc_dxt1_ext                     = int(0x8C4C)
	gl_compressed_srgb_s3tc_dxt1_nv                      = int(0x8C4C)
	gl_compressed_srgb_alpha_s3tc_dxt1_ext               = int(0x8C4D)
	gl_compressed_srgb_alpha_s3tc_dxt1_nv                = int(0x8C4D)
	gl_compressed_srgb_alpha_s3tc_dxt3_ext               = int(0x8C4E)
	gl_compressed_srgb_alpha_s3tc_dxt3_nv                = int(0x8C4E)
	gl_compressed_srgb_alpha_s3tc_dxt5_ext               = int(0x8C4F)
	gl_compressed_srgb_alpha_s3tc_dxt5_nv                = int(0x8C4F)
	gl_compressed_luminance_latc1_ext                    = int(0x8C70)
	gl_compressed_signed_luminance_latc1_ext             = int(0x8C71)
	gl_compressed_luminance_alpha_latc2_ext              = int(0x8C72)
	gl_compressed_signed_luminance_alpha_latc2_ext       = int(0x8C73)
	gl_tess_control_program_parameter_buffer_nv          = int(0x8C74)
	gl_tess_evaluation_program_parameter_buffer_nv       = int(0x8C75)
	gl_transform_feedback_varying_max_length             = int(0x8C76)
	gl_transform_feedback_varying_max_length_ext         = int(0x8C76)
	gl_back_primary_color_nv                             = int(0x8C77)
	gl_back_secondary_color_nv                           = int(0x8C78)
	gl_texture_coord_nv                                  = int(0x8C79)
	gl_clip_distance_nv                                  = int(0x8C7A)
	gl_vertex_id_nv                                      = int(0x8C7B)
	gl_primitive_id_nv                                   = int(0x8C7C)
	gl_generic_attrib_nv                                 = int(0x8C7D)
	gl_transform_feedback_attribs_nv                     = int(0x8C7E)
	gl_transform_feedback_buffer_mode                    = int(0x8C7F)
	gl_transform_feedback_buffer_mode_ext                = int(0x8C7F)
	gl_transform_feedback_buffer_mode_nv                 = int(0x8C7F)
	gl_max_transform_feedback_separate_components        = int(0x8C80)
	gl_max_transform_feedback_separate_components_ext    = int(0x8C80)
	gl_max_transform_feedback_separate_components_nv     = int(0x8C80)
	gl_active_varyings_nv                                = int(0x8C81)
	gl_active_varying_max_length_nv                      = int(0x8C82)
	gl_transform_feedback_varyings                       = int(0x8C83)
	gl_transform_feedback_varyings_ext                   = int(0x8C83)
	gl_transform_feedback_varyings_nv                    = int(0x8C83)
	gl_transform_feedback_buffer_start                   = int(0x8C84)
	gl_transform_feedback_buffer_start_ext               = int(0x8C84)
	gl_transform_feedback_buffer_start_nv                = int(0x8C84)
	gl_transform_feedback_buffer_size                    = int(0x8C85)
	gl_transform_feedback_buffer_size_ext                = int(0x8C85)
	gl_transform_feedback_buffer_size_nv                 = int(0x8C85)
	gl_transform_feedback_record_nv                      = int(0x8C86)
	gl_primitives_generated                              = int(0x8C87)
	gl_primitives_generated_ext                          = int(0x8C87)
	gl_primitives_generated_nv                           = int(0x8C87)
	gl_primitives_generated_oes                          = int(0x8C87)
	gl_transform_feedback_primitives_written             = int(0x8C88)
	gl_transform_feedback_primitives_written_ext         = int(0x8C88)
	gl_transform_feedback_primitives_written_nv          = int(0x8C88)
	gl_rasterizer_discard                                = int(0x8C89)
	gl_rasterizer_discard_ext                            = int(0x8C89)
	gl_rasterizer_discard_nv                             = int(0x8C89)
	gl_max_transform_feedback_interleaved_components     = int(0x8C8A)
	gl_max_transform_feedback_interleaved_components_ext = int(0x8C8A)
	gl_max_transform_feedback_interleaved_components_nv  = int(0x8C8A)
	gl_max_transform_feedback_separate_attribs           = int(0x8C8B)
	gl_max_transform_feedback_separate_attribs_ext       = int(0x8C8B)
	gl_max_transform_feedback_separate_attribs_nv        = int(0x8C8B)
	gl_interleaved_attribs                               = int(0x8C8C)
	gl_interleaved_attribs_ext                           = int(0x8C8C)
	gl_interleaved_attribs_nv                            = int(0x8C8C)
	gl_separate_attribs                                  = int(0x8C8D)
	gl_separate_attribs_ext                              = int(0x8C8D)
	gl_separate_attribs_nv                               = int(0x8C8D)
	gl_transform_feedback_buffer                         = int(0x8C8E)
	gl_transform_feedback_buffer_ext                     = int(0x8C8E)
	gl_transform_feedback_buffer_nv                      = int(0x8C8E)
	gl_transform_feedback_buffer_binding                 = int(0x8C8F)
	gl_transform_feedback_buffer_binding_ext             = int(0x8C8F)
	gl_transform_feedback_buffer_binding_nv              = int(0x8C8F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8C90" end="0x8C9F" vendor="QCOM" comment="For Affie Munshi. Reassigned from AMD to QCOM (bug 5874)" |>
pub const (
	gl_motion_estimation_search_block_x_qcom = int(0x8C90)
	gl_motion_estimation_search_block_y_qcom = int(0x8C91)
	gl_atc_rgb_amd                           = int(0x8C92)
	gl_atc_rgba_explicit_alpha_amd           = int(0x8C93)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8CA0" end="0x8CAF" vendor="ARB" |>
pub const (
	gl_point_sprite_coord_origin        = int(0x8CA0)
	gl_lower_left                       = int(0x8CA1)
	gl_lower_left_ext                   = int(0x8CA1)
	gl_upper_left                       = int(0x8CA2)
	gl_upper_left_ext                   = int(0x8CA2)
	gl_stencil_back_ref                 = int(0x8CA3)
	gl_stencil_back_value_mask          = int(0x8CA4)
	gl_stencil_back_writemask           = int(0x8CA5)
	gl_draw_framebuffer_binding         = int(0x8CA6)
	gl_draw_framebuffer_binding_angle   = int(0x8CA6)
	gl_draw_framebuffer_binding_apple   = int(0x8CA6)
	gl_draw_framebuffer_binding_ext     = int(0x8CA6)
	gl_draw_framebuffer_binding_nv      = int(0x8CA6)
	gl_framebuffer_binding              = int(0x8CA6)
	gl_framebuffer_binding_angle        = int(0x8CA6)
	gl_framebuffer_binding_ext          = int(0x8CA6)
	gl_framebuffer_binding_oes          = int(0x8CA6)
	gl_renderbuffer_binding             = int(0x8CA7)
	gl_renderbuffer_binding_angle       = int(0x8CA7)
	gl_renderbuffer_binding_ext         = int(0x8CA7)
	gl_renderbuffer_binding_oes         = int(0x8CA7)
	gl_read_framebuffer                 = int(0x8CA8)
	gl_read_framebuffer_angle           = int(0x8CA8)
	gl_read_framebuffer_apple           = int(0x8CA8)
	gl_read_framebuffer_ext             = int(0x8CA8)
	gl_read_framebuffer_nv              = int(0x8CA8)
	gl_draw_framebuffer                 = int(0x8CA9)
	gl_draw_framebuffer_angle           = int(0x8CA9)
	gl_draw_framebuffer_apple           = int(0x8CA9)
	gl_draw_framebuffer_ext             = int(0x8CA9)
	gl_draw_framebuffer_nv              = int(0x8CA9)
	gl_read_framebuffer_binding         = int(0x8CAA)
	gl_read_framebuffer_binding_angle   = int(0x8CAA)
	gl_read_framebuffer_binding_apple   = int(0x8CAA)
	gl_read_framebuffer_binding_ext     = int(0x8CAA)
	gl_read_framebuffer_binding_nv      = int(0x8CAA)
	gl_renderbuffer_coverage_samples_nv = int(0x8CAB)
	gl_renderbuffer_samples             = int(0x8CAB)
	gl_renderbuffer_samples_angle       = int(0x8CAB)
	gl_renderbuffer_samples_apple       = int(0x8CAB)
	gl_renderbuffer_samples_ext         = int(0x8CAB)
	gl_renderbuffer_samples_nv          = int(0x8CAB)
	gl_depth_component32f               = int(0x8CAC)
	gl_depth32f_stencil8                = int(0x8CAD)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8CD0" end="0x8D5F" vendor="ARB" comment="Framebuffer object specification + headroom" |>
pub const (
	gl_framebuffer_attachment_object_type               = int(0x8CD0)
	gl_framebuffer_attachment_object_type_ext           = int(0x8CD0)
	gl_framebuffer_attachment_object_type_oes           = int(0x8CD0)
	gl_framebuffer_attachment_object_name               = int(0x8CD1)
	gl_framebuffer_attachment_object_name_ext           = int(0x8CD1)
	gl_framebuffer_attachment_object_name_oes           = int(0x8CD1)
	gl_framebuffer_attachment_texture_level             = int(0x8CD2)
	gl_framebuffer_attachment_texture_level_ext         = int(0x8CD2)
	gl_framebuffer_attachment_texture_level_oes         = int(0x8CD2)
	gl_framebuffer_attachment_texture_cube_map_face     = int(0x8CD3)
	gl_framebuffer_attachment_texture_cube_map_face_ext = int(0x8CD3)
	gl_framebuffer_attachment_texture_cube_map_face_oes = int(0x8CD3)
	gl_framebuffer_attachment_texture_3d_zoffset_ext    = int(0x8CD4)
	gl_framebuffer_attachment_texture_3d_zoffset_oes    = int(0x8CD4)
	gl_framebuffer_attachment_texture_layer             = int(0x8CD4)
	gl_framebuffer_attachment_texture_layer_ext         = int(0x8CD4)
	gl_framebuffer_complete                             = int(0x8CD5)
	gl_framebuffer_complete_ext                         = int(0x8CD5)
	gl_framebuffer_complete_oes                         = int(0x8CD5)
	gl_framebuffer_incomplete_attachment                = int(0x8CD6)
	gl_framebuffer_incomplete_attachment_ext            = int(0x8CD6)
	gl_framebuffer_incomplete_attachment_oes            = int(0x8CD6)
	gl_framebuffer_incomplete_missing_attachment        = int(0x8CD7)
	gl_framebuffer_incomplete_missing_attachment_ext    = int(0x8CD7)
	gl_framebuffer_incomplete_missing_attachment_oes    = int(0x8CD7)
	gl_framebuffer_incomplete_dimensions                = int(0x8CD9)
	gl_framebuffer_incomplete_dimensions_ext            = int(0x8CD9)
	gl_framebuffer_incomplete_dimensions_oes            = int(0x8CD9)
	gl_framebuffer_incomplete_formats_ext               = int(0x8CDA)
	gl_framebuffer_incomplete_formats_oes               = int(0x8CDA)
	gl_framebuffer_incomplete_draw_buffer               = int(0x8CDB)
	gl_framebuffer_incomplete_draw_buffer_ext           = int(0x8CDB)
	gl_framebuffer_incomplete_draw_buffer_oes           = int(0x8CDB)
	gl_framebuffer_incomplete_read_buffer               = int(0x8CDC)
	gl_framebuffer_incomplete_read_buffer_ext           = int(0x8CDC)
	gl_framebuffer_incomplete_read_buffer_oes           = int(0x8CDC)
	gl_framebuffer_unsupported                          = int(0x8CDD)
	gl_framebuffer_unsupported_ext                      = int(0x8CDD)
	gl_framebuffer_unsupported_oes                      = int(0x8CDD)
	gl_max_color_attachments                            = int(0x8CDF)
	gl_max_color_attachments_ext                        = int(0x8CDF)
	gl_max_color_attachments_nv                         = int(0x8CDF)
	gl_color_attachment0                                = int(0x8CE0)
	gl_color_attachment0_ext                            = int(0x8CE0)
	gl_color_attachment0_nv                             = int(0x8CE0)
	gl_color_attachment0_oes                            = int(0x8CE0)
	gl_color_attachment1                                = int(0x8CE1)
	gl_color_attachment1_ext                            = int(0x8CE1)
	gl_color_attachment1_nv                             = int(0x8CE1)
	gl_color_attachment2                                = int(0x8CE2)
	gl_color_attachment2_ext                            = int(0x8CE2)
	gl_color_attachment2_nv                             = int(0x8CE2)
	gl_color_attachment3                                = int(0x8CE3)
	gl_color_attachment3_ext                            = int(0x8CE3)
	gl_color_attachment3_nv                             = int(0x8CE3)
	gl_color_attachment4                                = int(0x8CE4)
	gl_color_attachment4_ext                            = int(0x8CE4)
	gl_color_attachment4_nv                             = int(0x8CE4)
	gl_color_attachment5                                = int(0x8CE5)
	gl_color_attachment5_ext                            = int(0x8CE5)
	gl_color_attachment5_nv                             = int(0x8CE5)
	gl_color_attachment6                                = int(0x8CE6)
	gl_color_attachment6_ext                            = int(0x8CE6)
	gl_color_attachment6_nv                             = int(0x8CE6)
	gl_color_attachment7                                = int(0x8CE7)
	gl_color_attachment7_ext                            = int(0x8CE7)
	gl_color_attachment7_nv                             = int(0x8CE7)
	gl_color_attachment8                                = int(0x8CE8)
	gl_color_attachment8_ext                            = int(0x8CE8)
	gl_color_attachment8_nv                             = int(0x8CE8)
	gl_color_attachment9                                = int(0x8CE9)
	gl_color_attachment9_ext                            = int(0x8CE9)
	gl_color_attachment9_nv                             = int(0x8CE9)
	gl_color_attachment10                               = int(0x8CEA)
	gl_color_attachment10_ext                           = int(0x8CEA)
	gl_color_attachment10_nv                            = int(0x8CEA)
	gl_color_attachment11                               = int(0x8CEB)
	gl_color_attachment11_ext                           = int(0x8CEB)
	gl_color_attachment11_nv                            = int(0x8CEB)
	gl_color_attachment12                               = int(0x8CEC)
	gl_color_attachment12_ext                           = int(0x8CEC)
	gl_color_attachment12_nv                            = int(0x8CEC)
	gl_color_attachment13                               = int(0x8CED)
	gl_color_attachment13_ext                           = int(0x8CED)
	gl_color_attachment13_nv                            = int(0x8CED)
	gl_color_attachment14                               = int(0x8CEE)
	gl_color_attachment14_ext                           = int(0x8CEE)
	gl_color_attachment14_nv                            = int(0x8CEE)
	gl_color_attachment15                               = int(0x8CEF)
	gl_color_attachment15_ext                           = int(0x8CEF)
	gl_color_attachment15_nv                            = int(0x8CEF)
	gl_color_attachment16                               = int(0x8CF0)
	gl_color_attachment17                               = int(0x8CF1)
	gl_color_attachment18                               = int(0x8CF2)
	gl_color_attachment19                               = int(0x8CF3)
	gl_color_attachment20                               = int(0x8CF4)
	gl_color_attachment21                               = int(0x8CF5)
	gl_color_attachment22                               = int(0x8CF6)
	gl_color_attachment23                               = int(0x8CF7)
	gl_color_attachment24                               = int(0x8CF8)
	gl_color_attachment25                               = int(0x8CF9)
	gl_color_attachment26                               = int(0x8CFA)
	gl_color_attachment27                               = int(0x8CFB)
	gl_color_attachment28                               = int(0x8CFC)
	gl_color_attachment29                               = int(0x8CFD)
	gl_color_attachment30                               = int(0x8CFE)
	gl_color_attachment31                               = int(0x8CFF)
	gl_depth_attachment                                 = int(0x8D00)
	gl_depth_attachment_ext                             = int(0x8D00)
	gl_depth_attachment_oes                             = int(0x8D00)
	gl_stencil_attachment                               = int(0x8D20)
	gl_stencil_attachment_ext                           = int(0x8D20)
	gl_stencil_attachment_oes                           = int(0x8D20)
	gl_framebuffer                                      = int(0x8D40)
	gl_framebuffer_ext                                  = int(0x8D40)
	gl_framebuffer_oes                                  = int(0x8D40)
	gl_renderbuffer                                     = int(0x8D41)
	gl_renderbuffer_ext                                 = int(0x8D41)
	gl_renderbuffer_oes                                 = int(0x8D41)
	gl_renderbuffer_width                               = int(0x8D42)
	gl_renderbuffer_width_ext                           = int(0x8D42)
	gl_renderbuffer_width_oes                           = int(0x8D42)
	gl_renderbuffer_height                              = int(0x8D43)
	gl_renderbuffer_height_ext                          = int(0x8D43)
	gl_renderbuffer_height_oes                          = int(0x8D43)
	gl_renderbuffer_internal_format                     = int(0x8D44)
	gl_renderbuffer_internal_format_ext                 = int(0x8D44)
	gl_renderbuffer_internal_format_oes                 = int(0x8D44)
	gl_stencil_index1                                   = int(0x8D46)
	gl_stencil_index1_ext                               = int(0x8D46)
	gl_stencil_index1_oes                               = int(0x8D46)
	gl_stencil_index4                                   = int(0x8D47)
	gl_stencil_index4_ext                               = int(0x8D47)
	gl_stencil_index4_oes                               = int(0x8D47)
	gl_stencil_index8                                   = int(0x8D48)
	gl_stencil_index8_ext                               = int(0x8D48)
	gl_stencil_index8_oes                               = int(0x8D48)
	gl_stencil_index16                                  = int(0x8D49)
	gl_stencil_index16_ext                              = int(0x8D49)
	gl_renderbuffer_red_size                            = int(0x8D50)
	gl_renderbuffer_red_size_ext                        = int(0x8D50)
	gl_renderbuffer_red_size_oes                        = int(0x8D50)
	gl_renderbuffer_green_size                          = int(0x8D51)
	gl_renderbuffer_green_size_ext                      = int(0x8D51)
	gl_renderbuffer_green_size_oes                      = int(0x8D51)
	gl_renderbuffer_blue_size                           = int(0x8D52)
	gl_renderbuffer_blue_size_ext                       = int(0x8D52)
	gl_renderbuffer_blue_size_oes                       = int(0x8D52)
	gl_renderbuffer_alpha_size                          = int(0x8D53)
	gl_renderbuffer_alpha_size_ext                      = int(0x8D53)
	gl_renderbuffer_alpha_size_oes                      = int(0x8D53)
	gl_renderbuffer_depth_size                          = int(0x8D54)
	gl_renderbuffer_depth_size_ext                      = int(0x8D54)
	gl_renderbuffer_depth_size_oes                      = int(0x8D54)
	gl_renderbuffer_stencil_size                        = int(0x8D55)
	gl_renderbuffer_stencil_size_ext                    = int(0x8D55)
	gl_renderbuffer_stencil_size_oes                    = int(0x8D55)
	gl_framebuffer_incomplete_multisample               = int(0x8D56)
	gl_framebuffer_incomplete_multisample_angle         = int(0x8D56)
	gl_framebuffer_incomplete_multisample_apple         = int(0x8D56)
	gl_framebuffer_incomplete_multisample_ext           = int(0x8D56)
	gl_framebuffer_incomplete_multisample_nv            = int(0x8D56)
	gl_max_samples                                      = int(0x8D57)
	gl_max_samples_angle                                = int(0x8D57)
	gl_max_samples_apple                                = int(0x8D57)
	gl_max_samples_ext                                  = int(0x8D57)
	gl_max_samples_nv                                   = int(0x8D57)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8D60" end="0x8D6F" vendor="OES" |>
pub const (
	gl_texture_gen_str_oes                        = int(0x8D60)
	gl_half_float_oes                             = int(0x8D61)
	gl_rgb565_oes                                 = int(0x8D62)
	gl_rgb565                                     = int(0x8D62)
	gl_etc1_rgb8_oes                              = int(0x8D64)
	gl_texture_external_oes                       = int(0x8D65)
	gl_sampler_external_oes                       = int(0x8D66)
	gl_texture_binding_external_oes               = int(0x8D67)
	gl_required_texture_image_units_oes           = int(0x8D68)
	gl_primitive_restart_fixed_index              = int(0x8D69)
	gl_any_samples_passed_conservative            = int(0x8D6A)
	gl_any_samples_passed_conservative_ext        = int(0x8D6A)
	gl_max_element_index                          = int(0x8D6B)
	gl_framebuffer_attachment_texture_samples_ext = int(0x8D6C)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8D70" end="0x8DEF" vendor="NV" comment="For Pat Brown 2005/10/13" |>
pub const (
	gl_rgba32ui                                 = int(0x8D70)
	gl_rgba32ui_ext                             = int(0x8D70)
	gl_rgb32ui                                  = int(0x8D71)
	gl_rgb32ui_ext                              = int(0x8D71)
	gl_alpha32ui_ext                            = int(0x8D72)
	gl_intensity32ui_ext                        = int(0x8D73)
	gl_luminance32ui_ext                        = int(0x8D74)
	gl_luminance_alpha32ui_ext                  = int(0x8D75)
	gl_rgba16ui                                 = int(0x8D76)
	gl_rgba16ui_ext                             = int(0x8D76)
	gl_rgb16ui                                  = int(0x8D77)
	gl_rgb16ui_ext                              = int(0x8D77)
	gl_alpha16ui_ext                            = int(0x8D78)
	gl_intensity16ui_ext                        = int(0x8D79)
	gl_luminance16ui_ext                        = int(0x8D7A)
	gl_luminance_alpha16ui_ext                  = int(0x8D7B)
	gl_rgba8ui                                  = int(0x8D7C)
	gl_rgba8ui_ext                              = int(0x8D7C)
	gl_rgb8ui                                   = int(0x8D7D)
	gl_rgb8ui_ext                               = int(0x8D7D)
	gl_alpha8ui_ext                             = int(0x8D7E)
	gl_intensity8ui_ext                         = int(0x8D7F)
	gl_luminance8ui_ext                         = int(0x8D80)
	gl_luminance_alpha8ui_ext                   = int(0x8D81)
	gl_rgba32i                                  = int(0x8D82)
	gl_rgba32i_ext                              = int(0x8D82)
	gl_rgb32i                                   = int(0x8D83)
	gl_rgb32i_ext                               = int(0x8D83)
	gl_alpha32i_ext                             = int(0x8D84)
	gl_intensity32i_ext                         = int(0x8D85)
	gl_luminance32i_ext                         = int(0x8D86)
	gl_luminance_alpha32i_ext                   = int(0x8D87)
	gl_rgba16i                                  = int(0x8D88)
	gl_rgba16i_ext                              = int(0x8D88)
	gl_rgb16i                                   = int(0x8D89)
	gl_rgb16i_ext                               = int(0x8D89)
	gl_alpha16i_ext                             = int(0x8D8A)
	gl_intensity16i_ext                         = int(0x8D8B)
	gl_luminance16i_ext                         = int(0x8D8C)
	gl_luminance_alpha16i_ext                   = int(0x8D8D)
	gl_rgba8i                                   = int(0x8D8E)
	gl_rgba8i_ext                               = int(0x8D8E)
	gl_rgb8i                                    = int(0x8D8F)
	gl_rgb8i_ext                                = int(0x8D8F)
	gl_alpha8i_ext                              = int(0x8D90)
	gl_intensity8i_ext                          = int(0x8D91)
	gl_luminance8i_ext                          = int(0x8D92)
	gl_luminance_alpha8i_ext                    = int(0x8D93)
	gl_red_integer                              = int(0x8D94)
	gl_red_integer_ext                          = int(0x8D94)
	gl_green_integer                            = int(0x8D95)
	gl_green_integer_ext                        = int(0x8D95)
	gl_blue_integer                             = int(0x8D96)
	gl_blue_integer_ext                         = int(0x8D96)
	gl_alpha_integer                            = int(0x8D97)
	gl_alpha_integer_ext                        = int(0x8D97)
	gl_rgb_integer                              = int(0x8D98)
	gl_rgb_integer_ext                          = int(0x8D98)
	gl_rgba_integer                             = int(0x8D99)
	gl_rgba_integer_ext                         = int(0x8D99)
	gl_bgr_integer                              = int(0x8D9A)
	gl_bgr_integer_ext                          = int(0x8D9A)
	gl_bgra_integer                             = int(0x8D9B)
	gl_bgra_integer_ext                         = int(0x8D9B)
	gl_luminance_integer_ext                    = int(0x8D9C)
	gl_luminance_alpha_integer_ext              = int(0x8D9D)
	gl_rgba_integer_mode_ext                    = int(0x8D9E)
	gl_int_2_10_10_10_rev                       = int(0x8D9F)
	gl_max_program_parameter_buffer_bindings_nv = int(0x8DA0)
	gl_max_program_parameter_buffer_size_nv     = int(0x8DA1)
	gl_vertex_program_parameter_buffer_nv       = int(0x8DA2)
	gl_geometry_program_parameter_buffer_nv     = int(0x8DA3)
	gl_fragment_program_parameter_buffer_nv     = int(0x8DA4)
	gl_max_program_generic_attribs_nv           = int(0x8DA5)
	gl_max_program_generic_results_nv           = int(0x8DA6)
	gl_framebuffer_attachment_layered           = int(0x8DA7)
	gl_framebuffer_attachment_layered_arb       = int(0x8DA7)
	gl_framebuffer_attachment_layered_ext       = int(0x8DA7)
	gl_framebuffer_attachment_layered_oes       = int(0x8DA7)
	gl_framebuffer_incomplete_layer_targets     = int(0x8DA8)
	gl_framebuffer_incomplete_layer_targets_arb = int(0x8DA8)
	gl_framebuffer_incomplete_layer_targets_ext = int(0x8DA8)
	gl_framebuffer_incomplete_layer_targets_oes = int(0x8DA8)
	gl_framebuffer_incomplete_layer_count_arb   = int(0x8DA9)
	gl_framebuffer_incomplete_layer_count_ext   = int(0x8DA9)
	gl_layer_nv                                 = int(0x8DAA)
	gl_depth_component32f_nv                    = int(0x8DAB)
	gl_depth32f_stencil8_nv                     = int(0x8DAC)
	gl_float_32_unsigned_int_24_8_rev           = int(0x8DAD)
	gl_float_32_unsigned_int_24_8_rev_nv        = int(0x8DAD)
	gl_shader_include_arb                       = int(0x8DAE)
	gl_depth_buffer_float_mode_nv               = int(0x8DAF)
	gl_framebuffer_srgb                         = int(0x8DB9)
	gl_framebuffer_srgb_ext                     = int(0x8DB9)
	gl_framebuffer_srgb_capable_ext             = int(0x8DBA)
	gl_compressed_red_rgtc1                     = int(0x8DBB)
	gl_compressed_red_rgtc1_ext                 = int(0x8DBB)
	gl_compressed_signed_red_rgtc1              = int(0x8DBC)
	gl_compressed_signed_red_rgtc1_ext          = int(0x8DBC)
	gl_compressed_red_green_rgtc2_ext           = int(0x8DBD)
	gl_compressed_rg_rgtc2                      = int(0x8DBD)
	gl_compressed_signed_red_green_rgtc2_ext    = int(0x8DBE)
	gl_compressed_signed_rg_rgtc2               = int(0x8DBE)
	gl_sampler_1d_array                         = int(0x8DC0)
	gl_sampler_1d_array_ext                     = int(0x8DC0)
	gl_sampler_2d_array                         = int(0x8DC1)
	gl_sampler_2d_array_ext                     = int(0x8DC1)
	gl_sampler_buffer                           = int(0x8DC2)
	gl_sampler_buffer_ext                       = int(0x8DC2)
	gl_sampler_buffer_oes                       = int(0x8DC2)
	gl_sampler_1d_array_shadow                  = int(0x8DC3)
	gl_sampler_1d_array_shadow_ext              = int(0x8DC3)
	gl_sampler_2d_array_shadow                  = int(0x8DC4)
	gl_sampler_2d_array_shadow_ext              = int(0x8DC4)
	gl_sampler_2d_array_shadow_nv               = int(0x8DC4)
	gl_sampler_cube_shadow                      = int(0x8DC5)
	gl_sampler_cube_shadow_ext                  = int(0x8DC5)
	gl_sampler_cube_shadow_nv                   = int(0x8DC5)
	gl_unsigned_int_vec2                        = int(0x8DC6)
	gl_unsigned_int_vec2_ext                    = int(0x8DC6)
	gl_unsigned_int_vec3                        = int(0x8DC7)
	gl_unsigned_int_vec3_ext                    = int(0x8DC7)
	gl_unsigned_int_vec4                        = int(0x8DC8)
	gl_unsigned_int_vec4_ext                    = int(0x8DC8)
	gl_int_sampler_1d                           = int(0x8DC9)
	gl_int_sampler_1d_ext                       = int(0x8DC9)
	gl_int_sampler_2d                           = int(0x8DCA)
	gl_int_sampler_2d_ext                       = int(0x8DCA)
	gl_int_sampler_3d                           = int(0x8DCB)
	gl_int_sampler_3d_ext                       = int(0x8DCB)
	gl_int_sampler_cube                         = int(0x8DCC)
	gl_int_sampler_cube_ext                     = int(0x8DCC)
	gl_int_sampler_2d_rect                      = int(0x8DCD)
	gl_int_sampler_2d_rect_ext                  = int(0x8DCD)
	gl_int_sampler_1d_array                     = int(0x8DCE)
	gl_int_sampler_1d_array_ext                 = int(0x8DCE)
	gl_int_sampler_2d_array                     = int(0x8DCF)
	gl_int_sampler_2d_array_ext                 = int(0x8DCF)
	gl_int_sampler_buffer                       = int(0x8DD0)
	gl_int_sampler_buffer_ext                   = int(0x8DD0)
	gl_int_sampler_buffer_oes                   = int(0x8DD0)
	gl_unsigned_int_sampler_1d                  = int(0x8DD1)
	gl_unsigned_int_sampler_1d_ext              = int(0x8DD1)
	gl_unsigned_int_sampler_2d                  = int(0x8DD2)
	gl_unsigned_int_sampler_2d_ext              = int(0x8DD2)
	gl_unsigned_int_sampler_3d                  = int(0x8DD3)
	gl_unsigned_int_sampler_3d_ext              = int(0x8DD3)
	gl_unsigned_int_sampler_cube                = int(0x8DD4)
	gl_unsigned_int_sampler_cube_ext            = int(0x8DD4)
	gl_unsigned_int_sampler_2d_rect             = int(0x8DD5)
	gl_unsigned_int_sampler_2d_rect_ext         = int(0x8DD5)
	gl_unsigned_int_sampler_1d_array            = int(0x8DD6)
	gl_unsigned_int_sampler_1d_array_ext        = int(0x8DD6)
	gl_unsigned_int_sampler_2d_array            = int(0x8DD7)
	gl_unsigned_int_sampler_2d_array_ext        = int(0x8DD7)
	gl_unsigned_int_sampler_buffer              = int(0x8DD8)
	gl_unsigned_int_sampler_buffer_ext          = int(0x8DD8)
	gl_unsigned_int_sampler_buffer_oes          = int(0x8DD8)
	gl_geometry_shader                          = int(0x8DD9)
	gl_geometry_shader_arb                      = int(0x8DD9)
	gl_geometry_shader_ext                      = int(0x8DD9)
	gl_geometry_shader_oes                      = int(0x8DD9)
	gl_geometry_vertices_out_arb                = int(0x8DDA)
	gl_geometry_vertices_out_ext                = int(0x8DDA)
	gl_geometry_input_type_arb                  = int(0x8DDB)
	gl_geometry_input_type_ext                  = int(0x8DDB)
	gl_geometry_output_type_arb                 = int(0x8DDC)
	gl_geometry_output_type_ext                 = int(0x8DDC)
	gl_max_geometry_varying_components_arb      = int(0x8DDD)
	gl_max_geometry_varying_components_ext      = int(0x8DDD)
	gl_max_vertex_varying_components_arb        = int(0x8DDE)
	gl_max_vertex_varying_components_ext        = int(0x8DDE)
	gl_max_geometry_uniform_components          = int(0x8DDF)
	gl_max_geometry_uniform_components_arb      = int(0x8DDF)
	gl_max_geometry_uniform_components_ext      = int(0x8DDF)
	gl_max_geometry_uniform_components_oes      = int(0x8DDF)
	gl_max_geometry_output_vertices             = int(0x8DE0)
	gl_max_geometry_output_vertices_arb         = int(0x8DE0)
	gl_max_geometry_output_vertices_ext         = int(0x8DE0)
	gl_max_geometry_output_vertices_oes         = int(0x8DE0)
	gl_max_geometry_total_output_components     = int(0x8DE1)
	gl_max_geometry_total_output_components_arb = int(0x8DE1)
	gl_max_geometry_total_output_components_ext = int(0x8DE1)
	gl_max_geometry_total_output_components_oes = int(0x8DE1)
	gl_max_vertex_bindable_uniforms_ext         = int(0x8DE2)
	gl_max_fragment_bindable_uniforms_ext       = int(0x8DE3)
	gl_max_geometry_bindable_uniforms_ext       = int(0x8DE4)
	gl_active_subroutines                       = int(0x8DE5)
	gl_active_subroutine_uniforms               = int(0x8DE6)
	gl_max_subroutines                          = int(0x8DE7)
	gl_max_subroutine_uniform_locations         = int(0x8DE8)
	gl_named_string_length_arb                  = int(0x8DE9)
	gl_named_string_type_arb                    = int(0x8DEA)
	gl_max_bindable_uniform_size_ext            = int(0x8DED)
	gl_uniform_buffer_ext                       = int(0x8DEE)
	gl_uniform_buffer_binding_ext               = int(0x8DEF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8DF0" end="0x8E0F" vendor="OES" |>
pub const (
	gl_low_float                    = int(0x8DF0)
	gl_medium_float                 = int(0x8DF1)
	gl_high_float                   = int(0x8DF2)
	gl_low_int                      = int(0x8DF3)
	gl_medium_int                   = int(0x8DF4)
	gl_high_int                     = int(0x8DF5)
	gl_unsigned_int_10_10_10_2_oes  = int(0x8DF6)
	gl_int_10_10_10_2_oes           = int(0x8DF7)
	gl_shader_binary_formats        = int(0x8DF8)
	gl_num_shader_binary_formats    = int(0x8DF9)
	gl_shader_compiler              = int(0x8DFA)
	gl_max_vertex_uniform_vectors   = int(0x8DFB)
	gl_max_varying_vectors          = int(0x8DFC)
	gl_max_fragment_uniform_vectors = int(0x8DFD)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8E10" end="0x8E8F" vendor="NV" comment="For Michael Gold 2006/08/07" |>
pub const (
	gl_renderbuffer_color_samples_nv                       = int(0x8E10)
	gl_max_multisample_coverage_modes_nv                   = int(0x8E11)
	gl_multisample_coverage_modes_nv                       = int(0x8E12)
	gl_query_wait                                          = int(0x8E13)
	gl_query_wait_nv                                       = int(0x8E13)
	gl_query_no_wait                                       = int(0x8E14)
	gl_query_no_wait_nv                                    = int(0x8E14)
	gl_query_by_region_wait                                = int(0x8E15)
	gl_query_by_region_wait_nv                             = int(0x8E15)
	gl_query_by_region_no_wait                             = int(0x8E16)
	gl_query_by_region_no_wait_nv                          = int(0x8E16)
	gl_query_wait_inverted                                 = int(0x8E17)
	gl_query_no_wait_inverted                              = int(0x8E18)
	gl_query_by_region_wait_inverted                       = int(0x8E19)
	gl_query_by_region_no_wait_inverted                    = int(0x8E1A)
	gl_polygon_offset_clamp                                = int(0x8E1B)
	gl_polygon_offset_clamp_ext                            = int(0x8E1B)
	gl_max_combined_tess_control_uniform_components        = int(0x8E1E)
	gl_max_combined_tess_control_uniform_components_ext    = int(0x8E1E)
	gl_max_combined_tess_control_uniform_components_oes    = int(0x8E1E)
	gl_max_combined_tess_evaluation_uniform_components     = int(0x8E1F)
	gl_max_combined_tess_evaluation_uniform_components_ext = int(0x8E1F)
	gl_max_combined_tess_evaluation_uniform_components_oes = int(0x8E1F)
	gl_color_samples_nv                                    = int(0x8E20)
	gl_transform_feedback                                  = int(0x8E22)
	gl_transform_feedback_nv                               = int(0x8E22)
	gl_transform_feedback_buffer_paused                    = int(0x8E23)
	gl_transform_feedback_paused                           = int(0x8E23)
	gl_transform_feedback_buffer_paused_nv                 = int(0x8E23)
	gl_transform_feedback_buffer_active                    = int(0x8E24)
	gl_transform_feedback_active                           = int(0x8E24)
	gl_transform_feedback_buffer_active_nv                 = int(0x8E24)
	gl_transform_feedback_binding                          = int(0x8E25)
	gl_transform_feedback_binding_nv                       = int(0x8E25)
	gl_frame_nv                                            = int(0x8E26)
	gl_fields_nv                                           = int(0x8E27)
	gl_current_time_nv                                     = int(0x8E28)
	gl_timestamp                                           = int(0x8E28)
	gl_timestamp_ext                                       = int(0x8E28)
	gl_num_fill_streams_nv                                 = int(0x8E29)
	gl_present_time_nv                                     = int(0x8E2A)
	gl_present_duration_nv                                 = int(0x8E2B)
	gl_depth_component16_nonlinear_nv                      = int(0x8E2C)
	gl_program_matrix_ext                                  = int(0x8E2D)
	gl_transpose_program_matrix_ext                        = int(0x8E2E)
	gl_program_matrix_stack_depth_ext                      = int(0x8E2F)
	gl_texture_swizzle_r                                   = int(0x8E42)
	gl_texture_swizzle_r_ext                               = int(0x8E42)
	gl_texture_swizzle_g                                   = int(0x8E43)
	gl_texture_swizzle_g_ext                               = int(0x8E43)
	gl_texture_swizzle_b                                   = int(0x8E44)
	gl_texture_swizzle_b_ext                               = int(0x8E44)
	gl_texture_swizzle_a                                   = int(0x8E45)
	gl_texture_swizzle_a_ext                               = int(0x8E45)
	gl_texture_swizzle_rgba                                = int(0x8E46)
	gl_texture_swizzle_rgba_ext                            = int(0x8E46)
	gl_active_subroutine_uniform_locations                 = int(0x8E47)
	gl_active_subroutine_max_length                        = int(0x8E48)
	gl_active_subroutine_uniform_max_length                = int(0x8E49)
	gl_num_compatible_subroutines                          = int(0x8E4A)
	gl_compatible_subroutines                              = int(0x8E4B)
	gl_quads_follow_provoking_vertex_convention            = int(0x8E4C)
	gl_quads_follow_provoking_vertex_convention_ext        = int(0x8E4C)
	gl_first_vertex_convention                             = int(0x8E4D)
	gl_first_vertex_convention_ext                         = int(0x8E4D)
	gl_first_vertex_convention_oes                         = int(0x8E4D)
	gl_last_vertex_convention                              = int(0x8E4E)
	gl_last_vertex_convention_ext                          = int(0x8E4E)
	gl_last_vertex_convention_oes                          = int(0x8E4E)
	gl_provoking_vertex                                    = int(0x8E4F)
	gl_provoking_vertex_ext                                = int(0x8E4F)
	gl_sample_position                                     = int(0x8E50)
	gl_sample_position_nv                                  = int(0x8E50)
	gl_sample_location_arb                                 = int(0x8E50)
	gl_sample_location_nv                                  = int(0x8E50)
	gl_sample_mask                                         = int(0x8E51)
	gl_sample_mask_nv                                      = int(0x8E51)
	gl_sample_mask_value                                   = int(0x8E52)
	gl_sample_mask_value_nv                                = int(0x8E52)
	gl_texture_binding_renderbuffer_nv                     = int(0x8E53)
	gl_texture_renderbuffer_data_store_binding_nv          = int(0x8E54)
	gl_texture_renderbuffer_nv                             = int(0x8E55)
	gl_sampler_renderbuffer_nv                             = int(0x8E56)
	gl_int_sampler_renderbuffer_nv                         = int(0x8E57)
	gl_unsigned_int_sampler_renderbuffer_nv                = int(0x8E58)
	gl_max_sample_mask_words                               = int(0x8E59)
	gl_max_sample_mask_words_nv                            = int(0x8E59)
	gl_max_geometry_program_invocations_nv                 = int(0x8E5A)
	gl_max_geometry_shader_invocations                     = int(0x8E5A)
	gl_max_geometry_shader_invocations_ext                 = int(0x8E5A)
	gl_max_geometry_shader_invocations_oes                 = int(0x8E5A)
	gl_min_fragment_interpolation_offset                   = int(0x8E5B)
	gl_min_fragment_interpolation_offset_oes               = int(0x8E5B)
	gl_min_fragment_interpolation_offset_nv                = int(0x8E5B)
	gl_max_fragment_interpolation_offset                   = int(0x8E5C)
	gl_max_fragment_interpolation_offset_oes               = int(0x8E5C)
	gl_max_fragment_interpolation_offset_nv                = int(0x8E5C)
	gl_fragment_interpolation_offset_bits                  = int(0x8E5D)
	gl_fragment_interpolation_offset_bits_oes              = int(0x8E5D)
	gl_fragment_program_interpolation_offset_bits_nv       = int(0x8E5D)
	gl_min_program_texture_gather_offset                   = int(0x8E5E)
	gl_min_program_texture_gather_offset_arb               = int(0x8E5E)
	gl_min_program_texture_gather_offset_nv                = int(0x8E5E)
	gl_max_program_texture_gather_offset                   = int(0x8E5F)
	gl_max_program_texture_gather_offset_arb               = int(0x8E5F)
	gl_max_program_texture_gather_offset_nv                = int(0x8E5F)
	gl_max_mesh_uniform_blocks_nv                          = int(0x8E60)
	gl_max_mesh_texture_image_units_nv                     = int(0x8E61)
	gl_max_mesh_image_uniforms_nv                          = int(0x8E62)
	gl_max_mesh_uniform_components_nv                      = int(0x8E63)
	gl_max_mesh_atomic_counter_buffers_nv                  = int(0x8E64)
	gl_max_mesh_atomic_counters_nv                         = int(0x8E65)
	gl_max_mesh_shader_storage_blocks_nv                   = int(0x8E66)
	gl_max_combined_mesh_uniform_components_nv             = int(0x8E67)
	gl_max_task_uniform_blocks_nv                          = int(0x8E68)
	gl_max_task_texture_image_units_nv                     = int(0x8E69)
	gl_max_task_image_uniforms_nv                          = int(0x8E6A)
	gl_max_task_uniform_components_nv                      = int(0x8E6B)
	gl_max_task_atomic_counter_buffers_nv                  = int(0x8E6C)
	gl_max_task_atomic_counters_nv                         = int(0x8E6D)
	gl_max_task_shader_storage_blocks_nv                   = int(0x8E6E)
	gl_max_combined_task_uniform_components_nv             = int(0x8E6F)
	gl_max_transform_feedback_buffers                      = int(0x8E70)
	gl_max_vertex_streams                                  = int(0x8E71)
	gl_patch_vertices                                      = int(0x8E72)
	gl_patch_vertices_ext                                  = int(0x8E72)
	gl_patch_vertices_oes                                  = int(0x8E72)
	gl_patch_default_inner_level                           = int(0x8E73)
	gl_patch_default_inner_level_ext                       = int(0x8E73)
	gl_patch_default_outer_level                           = int(0x8E74)
	gl_patch_default_outer_level_ext                       = int(0x8E74)
	gl_tess_control_output_vertices                        = int(0x8E75)
	gl_tess_control_output_vertices_ext                    = int(0x8E75)
	gl_tess_control_output_vertices_oes                    = int(0x8E75)
	gl_tess_gen_mode                                       = int(0x8E76)
	gl_tess_gen_mode_ext                                   = int(0x8E76)
	gl_tess_gen_mode_oes                                   = int(0x8E76)
	gl_tess_gen_spacing                                    = int(0x8E77)
	gl_tess_gen_spacing_ext                                = int(0x8E77)
	gl_tess_gen_spacing_oes                                = int(0x8E77)
	gl_tess_gen_vertex_order                               = int(0x8E78)
	gl_tess_gen_vertex_order_ext                           = int(0x8E78)
	gl_tess_gen_vertex_order_oes                           = int(0x8E78)
	gl_tess_gen_point_mode                                 = int(0x8E79)
	gl_tess_gen_point_mode_ext                             = int(0x8E79)
	gl_tess_gen_point_mode_oes                             = int(0x8E79)
	gl_isolines                                            = int(0x8E7A)
	gl_isolines_ext                                        = int(0x8E7A)
	gl_isolines_oes                                        = int(0x8E7A)
	gl_fractional_odd                                      = int(0x8E7B)
	gl_fractional_odd_ext                                  = int(0x8E7B)
	gl_fractional_odd_oes                                  = int(0x8E7B)
	gl_fractional_even                                     = int(0x8E7C)
	gl_fractional_even_ext                                 = int(0x8E7C)
	gl_fractional_even_oes                                 = int(0x8E7C)
	gl_max_patch_vertices                                  = int(0x8E7D)
	gl_max_patch_vertices_ext                              = int(0x8E7D)
	gl_max_patch_vertices_oes                              = int(0x8E7D)
	gl_max_tess_gen_level                                  = int(0x8E7E)
	gl_max_tess_gen_level_ext                              = int(0x8E7E)
	gl_max_tess_gen_level_oes                              = int(0x8E7E)
	gl_max_tess_control_uniform_components                 = int(0x8E7F)
	gl_max_tess_control_uniform_components_ext             = int(0x8E7F)
	gl_max_tess_control_uniform_components_oes             = int(0x8E7F)
	gl_max_tess_evaluation_uniform_components              = int(0x8E80)
	gl_max_tess_evaluation_uniform_components_ext          = int(0x8E80)
	gl_max_tess_evaluation_uniform_components_oes          = int(0x8E80)
	gl_max_tess_control_texture_image_units                = int(0x8E81)
	gl_max_tess_control_texture_image_units_ext            = int(0x8E81)
	gl_max_tess_control_texture_image_units_oes            = int(0x8E81)
	gl_max_tess_evaluation_texture_image_units             = int(0x8E82)
	gl_max_tess_evaluation_texture_image_units_ext         = int(0x8E82)
	gl_max_tess_evaluation_texture_image_units_oes         = int(0x8E82)
	gl_max_tess_control_output_components                  = int(0x8E83)
	gl_max_tess_control_output_components_ext              = int(0x8E83)
	gl_max_tess_control_output_components_oes              = int(0x8E83)
	gl_max_tess_patch_components                           = int(0x8E84)
	gl_max_tess_patch_components_ext                       = int(0x8E84)
	gl_max_tess_patch_components_oes                       = int(0x8E84)
	gl_max_tess_control_total_output_components            = int(0x8E85)
	gl_max_tess_control_total_output_components_ext        = int(0x8E85)
	gl_max_tess_control_total_output_components_oes        = int(0x8E85)
	gl_max_tess_evaluation_output_components               = int(0x8E86)
	gl_max_tess_evaluation_output_components_ext           = int(0x8E86)
	gl_max_tess_evaluation_output_components_oes           = int(0x8E86)
	gl_tess_evaluation_shader                              = int(0x8E87)
	gl_tess_evaluation_shader_ext                          = int(0x8E87)
	gl_tess_evaluation_shader_oes                          = int(0x8E87)
	gl_tess_control_shader                                 = int(0x8E88)
	gl_tess_control_shader_ext                             = int(0x8E88)
	gl_tess_control_shader_oes                             = int(0x8E88)
	gl_max_tess_control_uniform_blocks                     = int(0x8E89)
	gl_max_tess_control_uniform_blocks_ext                 = int(0x8E89)
	gl_max_tess_control_uniform_blocks_oes                 = int(0x8E89)
	gl_max_tess_evaluation_uniform_blocks                  = int(0x8E8A)
	gl_max_tess_evaluation_uniform_blocks_ext              = int(0x8E8A)
	gl_max_tess_evaluation_uniform_blocks_oes              = int(0x8E8A)
	gl_compressed_rgba_bptc_unorm                          = int(0x8E8C)
	gl_compressed_rgba_bptc_unorm_arb                      = int(0x8E8C)
	gl_compressed_rgba_bptc_unorm_ext                      = int(0x8E8C)
	gl_compressed_srgb_alpha_bptc_unorm                    = int(0x8E8D)
	gl_compressed_srgb_alpha_bptc_unorm_arb                = int(0x8E8D)
	gl_compressed_srgb_alpha_bptc_unorm_ext                = int(0x8E8D)
	gl_compressed_rgb_bptc_signed_float                    = int(0x8E8E)
	gl_compressed_rgb_bptc_signed_float_arb                = int(0x8E8E)
	gl_compressed_rgb_bptc_signed_float_ext                = int(0x8E8E)
	gl_compressed_rgb_bptc_unsigned_float                  = int(0x8E8F)
	gl_compressed_rgb_bptc_unsigned_float_arb              = int(0x8E8F)
	gl_compressed_rgb_bptc_unsigned_float_ext              = int(0x8E8F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8EA0" end="0x8EAF" vendor="IMG" |>
pub const (
	gl_trp_img                      = int(0x8EA0)
	gl_trp_error_context_reset_img  = int(0x8EA1)
	gl_trp_unsupported_context_img  = int(0x8EA2)
	gl_pvric_signature_mismatch_img = int(0x8EA3)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8ED0" end="0x8F4F" vendor="NV" comment="For Pat Brown, Khronos bug 3191" |>
pub const (
	gl_coverage_component_nv                             = int(0x8ED0)
	gl_coverage_component4_nv                            = int(0x8ED1)
	gl_coverage_attachment_nv                            = int(0x8ED2)
	gl_coverage_buffers_nv                               = int(0x8ED3)
	gl_coverage_samples_nv                               = int(0x8ED4)
	gl_coverage_all_fragments_nv                         = int(0x8ED5)
	gl_coverage_edge_fragments_nv                        = int(0x8ED6)
	gl_coverage_automatic_nv                             = int(0x8ED7)
	gl_inclusive_ext                                     = int(0x8F10)
	gl_exclusive_ext                                     = int(0x8F11)
	gl_window_rectangle_ext                              = int(0x8F12)
	gl_window_rectangle_mode_ext                         = int(0x8F13)
	gl_max_window_rectangles_ext                         = int(0x8F14)
	gl_num_window_rectangles_ext                         = int(0x8F15)
	gl_buffer_gpu_address_nv                             = int(0x8F1D)
	gl_vertex_attrib_array_unified_nv                    = int(0x8F1E)
	gl_element_array_unified_nv                          = int(0x8F1F)
	gl_vertex_attrib_array_address_nv                    = int(0x8F20)
	gl_vertex_array_address_nv                           = int(0x8F21)
	gl_normal_array_address_nv                           = int(0x8F22)
	gl_color_array_address_nv                            = int(0x8F23)
	gl_index_array_address_nv                            = int(0x8F24)
	gl_texture_coord_array_address_nv                    = int(0x8F25)
	gl_edge_flag_array_address_nv                        = int(0x8F26)
	gl_secondary_color_array_address_nv                  = int(0x8F27)
	gl_fog_coord_array_address_nv                        = int(0x8F28)
	gl_element_array_address_nv                          = int(0x8F29)
	gl_vertex_attrib_array_length_nv                     = int(0x8F2A)
	gl_vertex_array_length_nv                            = int(0x8F2B)
	gl_normal_array_length_nv                            = int(0x8F2C)
	gl_color_array_length_nv                             = int(0x8F2D)
	gl_index_array_length_nv                             = int(0x8F2E)
	gl_texture_coord_array_length_nv                     = int(0x8F2F)
	gl_edge_flag_array_length_nv                         = int(0x8F30)
	gl_secondary_color_array_length_nv                   = int(0x8F31)
	gl_fog_coord_array_length_nv                         = int(0x8F32)
	gl_element_array_length_nv                           = int(0x8F33)
	gl_gpu_address_nv                                    = int(0x8F34)
	gl_max_shader_buffer_address_nv                      = int(0x8F35)
	gl_copy_read_buffer                                  = int(0x8F36)
	gl_copy_read_buffer_nv                               = int(0x8F36)
	gl_copy_read_buffer_binding                          = int(0x8F36)
	gl_copy_write_buffer                                 = int(0x8F37)
	gl_copy_write_buffer_nv                              = int(0x8F37)
	gl_copy_write_buffer_binding                         = int(0x8F37)
	gl_max_image_units                                   = int(0x8F38)
	gl_max_image_units_ext                               = int(0x8F38)
	gl_max_combined_image_units_and_fragment_outputs     = int(0x8F39)
	gl_max_combined_image_units_and_fragment_outputs_ext = int(0x8F39)
	gl_max_combined_shader_output_resources              = int(0x8F39)
	gl_image_binding_name                                = int(0x8F3A)
	gl_image_binding_name_ext                            = int(0x8F3A)
	gl_image_binding_level                               = int(0x8F3B)
	gl_image_binding_level_ext                           = int(0x8F3B)
	gl_image_binding_layered                             = int(0x8F3C)
	gl_image_binding_layered_ext                         = int(0x8F3C)
	gl_image_binding_layer                               = int(0x8F3D)
	gl_image_binding_layer_ext                           = int(0x8F3D)
	gl_image_binding_access                              = int(0x8F3E)
	gl_image_binding_access_ext                          = int(0x8F3E)
	gl_draw_indirect_buffer                              = int(0x8F3F)
	gl_draw_indirect_unified_nv                          = int(0x8F40)
	gl_draw_indirect_address_nv                          = int(0x8F41)
	gl_draw_indirect_length_nv                           = int(0x8F42)
	gl_draw_indirect_buffer_binding                      = int(0x8F43)
	gl_max_program_subroutine_parameters_nv              = int(0x8F44)
	gl_max_program_subroutine_num_nv                     = int(0x8F45)
	gl_double_mat2                                       = int(0x8F46)
	gl_double_mat2_ext                                   = int(0x8F46)
	gl_double_mat3                                       = int(0x8F47)
	gl_double_mat3_ext                                   = int(0x8F47)
	gl_double_mat4                                       = int(0x8F48)
	gl_double_mat4_ext                                   = int(0x8F48)
	gl_double_mat2x3                                     = int(0x8F49)
	gl_double_mat2x3_ext                                 = int(0x8F49)
	gl_double_mat2x4                                     = int(0x8F4A)
	gl_double_mat2x4_ext                                 = int(0x8F4A)
	gl_double_mat3x2                                     = int(0x8F4B)
	gl_double_mat3x2_ext                                 = int(0x8F4B)
	gl_double_mat3x4                                     = int(0x8F4C)
	gl_double_mat3x4_ext                                 = int(0x8F4C)
	gl_double_mat4x2                                     = int(0x8F4D)
	gl_double_mat4x2_ext                                 = int(0x8F4D)
	gl_double_mat4x3                                     = int(0x8F4E)
	gl_double_mat4x3_ext                                 = int(0x8F4E)
	gl_vertex_binding_buffer                             = int(0x8F4F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8F60" end="0x8F6F" vendor="ARM" comment="For Remi Pedersen, Khronos bug 3745" |>
pub const (
	gl_mali_shader_binary_arm                                    = int(0x8F60)
	gl_mali_program_binary_arm                                   = int(0x8F61)
	gl_max_shader_pixel_local_storage_fast_size_ext              = int(0x8F63)
	gl_shader_pixel_local_storage_ext                            = int(0x8F64)
	gl_fetch_per_sample_arm                                      = int(0x8F65)
	gl_fragment_shader_framebuffer_fetch_mrt_arm                 = int(0x8F66)
	gl_max_shader_pixel_local_storage_size_ext                   = int(0x8F67)
	gl_texture_astc_decode_precision_ext                         = int(0x8F69)
	gl_texture_unnormalized_coordinates_arm                      = int(0x8F6A)
	gl_num_surface_compression_fixed_rates_ext                   = int(0x8F6E)
	gl_fragment_shading_rate_non_trivial_combiners_supported_ext = int(0x8F6F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8F90" end="0x8F9F" vendor="ARB" |>
pub const (
	gl_red_snorm                                 = int(0x8F90)
	gl_rg_snorm                                  = int(0x8F91)
	gl_rgb_snorm                                 = int(0x8F92)
	gl_rgba_snorm                                = int(0x8F93)
	gl_r8_snorm                                  = int(0x8F94)
	gl_rg8_snorm                                 = int(0x8F95)
	gl_rgb8_snorm                                = int(0x8F96)
	gl_rgba8_snorm                               = int(0x8F97)
	gl_r16_snorm                                 = int(0x8F98)
	gl_r16_snorm_ext                             = int(0x8F98)
	gl_rg16_snorm                                = int(0x8F99)
	gl_rg16_snorm_ext                            = int(0x8F99)
	gl_rgb16_snorm                               = int(0x8F9A)
	gl_rgb16_snorm_ext                           = int(0x8F9A)
	gl_rgba16_snorm                              = int(0x8F9B)
	gl_rgba16_snorm_ext                          = int(0x8F9B)
	gl_signed_normalized                         = int(0x8F9C)
	gl_primitive_restart                         = int(0x8F9D)
	gl_primitive_restart_index                   = int(0x8F9E)
	gl_max_program_texture_gather_components_arb = int(0x8F9F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8FA0" end="0x8FBF" vendor="QCOM" comment="For Maurice Ribble, bug 4512" |>
pub const (
	gl_perfmon_global_mode_qcom               = int(0x8FA0)
	gl_max_shader_subsampled_image_units_qcom = int(0x8FA1)
	gl_binning_control_hint_qcom              = int(0x8FB0)
	gl_cpu_optimized_qcom                     = int(0x8FB1)
	gl_gpu_optimized_qcom                     = int(0x8FB2)
	gl_render_direct_to_framebuffer_qcom      = int(0x8FB3)
	gl_gpu_disjoint_ext                       = int(0x8FBB)
	gl_sr8_ext                                = int(0x8FBD)
	gl_srg8_ext                               = int(0x8FBE)
	gl_texture_format_srgb_override_ext       = int(0x8FBF)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8FC0" end="0x8FDF" vendor="VIV" comment="For Frido Garritsen, bug 4526" |>
pub const (
	gl_shader_binary_viv = int(0x8FC4)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x8FE0" end="0x8FFF" vendor="NV" comment="For Pat Brown, bug 4935" |>
pub const (
	gl_int8_nv                 = int(0x8FE0)
	gl_int8_vec2_nv            = int(0x8FE1)
	gl_int8_vec3_nv            = int(0x8FE2)
	gl_int8_vec4_nv            = int(0x8FE3)
	gl_int16_nv                = int(0x8FE4)
	gl_int16_vec2_nv           = int(0x8FE5)
	gl_int16_vec3_nv           = int(0x8FE6)
	gl_int16_vec4_nv           = int(0x8FE7)
	gl_int64_vec2_arb          = int(0x8FE9)
	gl_int64_vec2_nv           = int(0x8FE9)
	gl_int64_vec3_arb          = int(0x8FEA)
	gl_int64_vec3_nv           = int(0x8FEA)
	gl_int64_vec4_arb          = int(0x8FEB)
	gl_int64_vec4_nv           = int(0x8FEB)
	gl_unsigned_int8_nv        = int(0x8FEC)
	gl_unsigned_int8_vec2_nv   = int(0x8FED)
	gl_unsigned_int8_vec3_nv   = int(0x8FEE)
	gl_unsigned_int8_vec4_nv   = int(0x8FEF)
	gl_unsigned_int16_nv       = int(0x8FF0)
	gl_unsigned_int16_vec2_nv  = int(0x8FF1)
	gl_unsigned_int16_vec3_nv  = int(0x8FF2)
	gl_unsigned_int16_vec4_nv  = int(0x8FF3)
	gl_unsigned_int64_vec2_arb = int(0x8FF5)
	gl_unsigned_int64_vec2_nv  = int(0x8FF5)
	gl_unsigned_int64_vec3_arb = int(0x8FF6)
	gl_unsigned_int64_vec3_nv  = int(0x8FF6)
	gl_unsigned_int64_vec4_arb = int(0x8FF7)
	gl_unsigned_int64_vec4_nv  = int(0x8FF7)
	gl_float16_nv              = int(0x8FF8)
	gl_float16_vec2_nv         = int(0x8FF9)
	gl_float16_vec3_nv         = int(0x8FFA)
	gl_float16_vec4_nv         = int(0x8FFB)
	gl_double_vec2             = int(0x8FFC)
	gl_double_vec2_ext         = int(0x8FFC)
	gl_double_vec3             = int(0x8FFD)
	gl_double_vec3_ext         = int(0x8FFD)
	gl_double_vec4             = int(0x8FFE)
	gl_double_vec4_ext         = int(0x8FFE)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x9000" end="0x901F" vendor="AMD" comment="For Bill Licea-Kane" |>
pub const (
	gl_sampler_buffer_amd                      = int(0x9001)
	gl_int_sampler_buffer_amd                  = int(0x9002)
	gl_unsigned_int_sampler_buffer_amd         = int(0x9003)
	gl_tessellation_mode_amd                   = int(0x9004)
	gl_tessellation_factor_amd                 = int(0x9005)
	gl_discrete_amd                            = int(0x9006)
	gl_continuous_amd                          = int(0x9007)
	gl_texture_cube_map_array                  = int(0x9009)
	gl_texture_cube_map_array_arb              = int(0x9009)
	gl_texture_cube_map_array_ext              = int(0x9009)
	gl_texture_cube_map_array_oes              = int(0x9009)
	gl_texture_binding_cube_map_array          = int(0x900A)
	gl_texture_binding_cube_map_array_arb      = int(0x900A)
	gl_texture_binding_cube_map_array_ext      = int(0x900A)
	gl_texture_binding_cube_map_array_oes      = int(0x900A)
	gl_proxy_texture_cube_map_array            = int(0x900B)
	gl_proxy_texture_cube_map_array_arb        = int(0x900B)
	gl_sampler_cube_map_array                  = int(0x900C)
	gl_sampler_cube_map_array_arb              = int(0x900C)
	gl_sampler_cube_map_array_ext              = int(0x900C)
	gl_sampler_cube_map_array_oes              = int(0x900C)
	gl_sampler_cube_map_array_shadow           = int(0x900D)
	gl_sampler_cube_map_array_shadow_arb       = int(0x900D)
	gl_sampler_cube_map_array_shadow_ext       = int(0x900D)
	gl_sampler_cube_map_array_shadow_oes       = int(0x900D)
	gl_int_sampler_cube_map_array              = int(0x900E)
	gl_int_sampler_cube_map_array_arb          = int(0x900E)
	gl_int_sampler_cube_map_array_ext          = int(0x900E)
	gl_int_sampler_cube_map_array_oes          = int(0x900E)
	gl_unsigned_int_sampler_cube_map_array     = int(0x900F)
	gl_unsigned_int_sampler_cube_map_array_arb = int(0x900F)
	gl_unsigned_int_sampler_cube_map_array_ext = int(0x900F)
	gl_unsigned_int_sampler_cube_map_array_oes = int(0x900F)
	gl_alpha_snorm                             = int(0x9010)
	gl_luminance_snorm                         = int(0x9011)
	gl_luminance_alpha_snorm                   = int(0x9012)
	gl_intensity_snorm                         = int(0x9013)
	gl_alpha8_snorm                            = int(0x9014)
	gl_luminance8_snorm                        = int(0x9015)
	gl_luminance8_alpha8_snorm                 = int(0x9016)
	gl_intensity8_snorm                        = int(0x9017)
	gl_alpha16_snorm                           = int(0x9018)
	gl_luminance16_snorm                       = int(0x9019)
	gl_luminance16_alpha16_snorm               = int(0x901A)
	gl_intensity16_snorm                       = int(0x901B)
	gl_factor_min_amd                          = int(0x901C)
	gl_factor_max_amd                          = int(0x901D)
	gl_depth_clamp_near_amd                    = int(0x901E)
	gl_depth_clamp_far_amd                     = int(0x901F)
)

// [ENUM SECTION (in V its just constants)] -> namespace="GL" start="0x9020" end="0x90FF" vendor="NV" comment="For Pat Brown, bug 4935" |>
pub const (
	gl_video_buffer_nv                              = int(0x9020)
	gl_video_buffer_binding_nv                      = int(0x9021)
	gl_field_upper_nv                               = int(0x9022)
	gl_field_lower_nv                               = int(0x9023)
	gl_num_video_capture_streams_nv                 = int(0x9024)
	gl_next_video_capture_buffer_status_nv          = int(0x9025)
	gl_video_capture_to_422_supported_nv            = int(0x9026)
	gl_last_video_capture_status_nv                 = int(0x9027)
	gl_video_buffer_pitch_nv                        = int(0x9028)
	gl_video_color_conversion_matrix_nv             = int(0x9029)
	gl_video_color_conversion_max_nv                = int(0x902A)
	gl_video_color_conversion_min_nv                = int(0x902B)
	gl_video_color_conversion_offset_nv             = int(0x902C)
	gl_video_buffer_internal_format_nv              = int(0x902D)
	gl_partial_success_nv                           = int(0x902E)
	gl_success_nv                                   = int(0x902F)
	gl_failure_nv                                   = int(0x9030)
	gl_ycbycr8_422_nv                               = int(0x9031)
	gl_ycbaycr8a_4224_nv                            = int(0x9032)
	gl_z6y10z6cb10z6y10z6cr10_422_nv                = int(0x9033)
	gl_z6y10z6cb10z6a10z6y10z6cr10z6a10_4224_nv     = int(0x9034)
	gl_z4y12z4cb12z4y12z4cr12_422_nv                = int(0x9035)
	gl_z4y12z4cb12z4a12z4y12z4cr12z4a12_4224_nv     = int(0x9036)
	gl_z4y12z4cb12z4cr12_444_nv                     = int(0x9037)
	gl_video_capture_frame_width_nv                 = int(0x9038)
	gl_video_capture_frame_height_nv                = int(0x9039)
	gl_video_capture_field_upper_height_nv          = int(0x903A)
	gl_video_capture_field_lower_height_nv          = int(0x903B)
	gl_video_capture_surface_origin_nv              = int(0x903C)
	gl_texture_coverage_samples_nv                  = int(0x9045)
	gl_texture_color_samples_nv                     = int(0x9046)
	gl_gpu_memory_info_dedicated_vidmem_nvx         = int(0x9047)
	gl_gpu_memory_info_total_available_memory_nvx   = int(0x9048)
	gl_gpu_memory_info_current_available_vidmem_nvx = int(0x9049)
	gl_gpu_memory_info_eviction_count_nvx           = int(0x904A)
	gl_gpu_memory_info_evicted_memory_nvx           = int(0x904B)
	gl_image_1d                                     = int(0x904C)
	gl_image_1d_ext                                 = int(0x904C)
	gl_image_2d                                     = int(0x904D)
	gl_image_2d_ext                                 = int(0x904D)
	gl_image_3d                                     = int(0x904E)
	gl_image_3d_ext                                 = int(0x904E)
	gl_image_2d_rect                                = int(0x904F)
	gl_image_2d_rect_ext                            = int(0x904F)
	gl_image_cube                                   = int(0x9050)
	gl_image_cube_ext                               = int(0x9050)
	gl_image_buffer                                 = int(0x9051)
	gl_image_buffer_ext                             = int(0x9051)
	gl_image_buffer_oes                             = int(0x9051)
	gl_image_1d_array                               = int(0x9052)
	gl_image_1d_array_ext                           = int(0x9052)
	gl_image_2d_array                               = int(0x9053)
	gl_image_2d_array_ext                           = int(0x9053)
	gl_image_cube_map_array                         = int(0x9054)
	gl_image_cube_map_array_ext                     = int(0x9054)
	gl_image_cube_map_array_oes                     = int(0x9054)
	gl_image_2d_multisample                         = int(0x9055)
	gl_image_2d_multisample_ext                     = int(0x9055)
	gl_image_2d_multisample_array                   = int(0x9056)
	gl_image_2d_multisample_array_ext               = int(0x9056)
	gl_int_image_1d                                 = int(0x9057)
	gl_int_image_1d_ext                             = int(0x9057)
	gl_int_image_2d                                 = int(0x9058)
	gl_int_image_2d_ext                             = int(0x9058)
	gl_int_image_3d                                 = int(0x9059)
	gl_int_image_3d_ext                             = int(0x9059)
	gl_int_image_2d_rect                            = int(0x905A)
	gl_int_image_2d_rect_ext                        = int(0x905A)
	gl_int_image_cube                               = int(0x905B)
	gl_int_image_cube_ext                           = int(0x905B)
	gl_int_image_buffer                             = int(0x905C)
	gl_int_image_buffer_ext                         = int(0x905C)
	gl_int_image_buffer_oes                         = int(0x905C)
	gl_int_image_1d_array                           = int(0x905D)
	gl_int_image_1d_array_ext                       = int(0x905D)
	gl_int_image_2d_array                           = int(0x905E)
	gl_int_image_2d_array_ext                       = int(0x905E)
	gl_int_image_cube_map_array                     = int(0x905F)
	gl_int_image_cube_map_array_ext                 = int(0x905F)
	gl_int_image_cube_map_array_oes                 = int(0x905F)
	gl_int_image_2d_multisample                     = int(0x9060)
	gl_int_image_2d_multisample_ext                 = int(0x9060)
	gl_int_image_2d_multisample_array               = int(0x9061)
	gl_int_image_2d_multisample_array_ext           = int(0x9061)
	gl_unsigned_int_image_1d                        = int(0x9062)
	gl_unsigned_int_image_1d_ext                    = int(0x9062)
	gl_unsigned_int_image_2d                        = int(0x9063)
	gl_unsigned_int_image_2d_ext                    = int(0x9063)
	gl_unsigned_int_image_3d                        = int(0x9064)
	gl_unsigned_int_image_3d_ext                    = int(0x9064)
	gl_unsigned_int_image_2d_rect                   = int(0x9065)
	gl_unsigned_int_image_2d_rect_ext               = int(0x9065)
	gl_unsigned_int_image_cube                      = int(0x9066)
	gl_unsigned_int_image_cube_ext                  = int(0x9066)
	gl_unsigned_int_image_buffer                    = int(0x9067)
	gl_unsigned_int_image_buffer_ext                = int(0x9067)
	gl_unsigned_int_image_buffer_oes                = int(0x9067)
	gl_unsigned_int_image_1d_array                  = int(0x9068)
	gl_unsigned_int_image_1d_array_ext              = int(0x9068)
	gl_unsigned_int_image_2d_array                  = int(0x9069)
	gl_unsigned_int_image_2d_array_ext              = int(0x9069)
	gl_unsigned_int_image_cube_map_array            = int(0x906A)
	gl_unsigned_int_image_cube_map_array_ext        = int(0x906A)
	gl_unsigned_int_image_cube_map_array_oes        = int(0x906A)
	gl_unsigned_int_image_2d_multisample            = int(0x906B)
	gl_unsigned_int_image_2d_multisample_ext        = int(0x906B)
	gl_unsigned_int_image_2d_multisample_array      = int(0x906C)
	gl_unsigned_int_image_2d_multisample_array_ext  = int(0x906C)
	gl_max_image_samples                            = int(0x906D)
	gl_max_image_samples_ext                        = int(0x906D)
	gl_image_binding_format                         = int(0x906E)
	gl_image_binding_format_ext                     = int(0x906E)
	gl_rgb10_a2ui                                   = int(0x906F)
	gl_path_format_svg_nv                           = int(0x9070)
	gl_path_format_ps_nv                            = int(0x9071)
	gl_standard_font_name_nv                        = int(0x9072)
	gl_system_font_name_nv                          = int(0x9073)
	gl_file_name_nv                                 = int(0x9074)
	gl_path_stroke_width_nv                         = int(0x9075)
	gl_path_end_caps_nv                             = int(0x9076)
	gl_path_initial_end_cap_nv                      = int(0x9077)
	gl_path_terminal_end_cap_nv                     = int(0x9078)
	gl_path_join_style_nv                           = int(0x9079)
	gl_path_miter_limit_nv                          = int(0x907A)
	gl_path_dash_caps_nv                            = int(0x907B)
	gl_path_initial_dash_cap_nv                     = int(0x907C)
	gl_path_terminal_dash_cap_nv                    = int(0x907D)
	gl_path_dash_offset_nv                          = int(0x907E)
	gl_path_client_length_nv                        = int(0x907F)
	gl_path_fill_mode_nv                            = int(0x9080)
	gl_path_fill_mask_nv                            = int(0x9081)
	gl_path_fill_cover_mode_nv                      = int(0x9082)
	gl_path_stroke_cover_mode_nv                    = int(0x9083)
)
