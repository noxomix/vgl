module vgl

#flag -I @VMODROOT/c/
#define GLAD_GL_IMPLEMENTATION
#include "/gl/gl.h"
#include "fallback.h"

#include <math.h>
#include <stdlib.h>
#include <stdio.h>
#include <string.h>
